Vim�UnDo� 8
A��ʭ�<(8���B7mt��$KQkm&��;   ?                                   ^X    _�                              ����                                                                                                                                                                                                                                                                                                                                                             ^W    �                (architecture Behavioral of split_1to8 is�                end split_1to8;�                entity split_1to8 is5��