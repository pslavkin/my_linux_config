Vim�UnDo� ��f[V�V��4=Ɵ�;�eWtc��X�=�ZP   F   #m_axis_config_tdata  <= "00000001";   C   "      N       N   N   N    ^-�(    _�                             ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �                )architecture Behavioral of join_8from2 is�                end join_8from2;�                entity join_8from2 is5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ^��    �          >      library IEEE;   use IEEE.STD_LOGIC_1164.ALL;5�_�                    +   @    ����                                                                                                                                                                                                                                                                                                                                                  V        ^��     �   *   ,   >      B                     bitCounter                 := bitCounter + 2;5�_�                    (   @    ����                                                                                                                                                                                                                                                                                                                                                  V        ^��     �   (   *   >    5�_�                    )        ����                                                                                                                                                                                                                                                                                                                                                  V        ^��     �   (   )           5�_�                       1    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �      	   >      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�                    )   "    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �   (   *   >    �   )   *   >    5�_�      	              )       ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �   (   *   ?      B                     bitCounter                 := bitCounter + 1;5�_�      
           	   )   #    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�#     �   (   *   ?      E                     if bitCounter                 := bitCounter + 1;5�_�   	              
   )   #    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�$     �   (   *   ?      '                     if bitCounter + 1;5�_�   
                 )   &    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�'     �   (   *   ?      '                     if bitCounter = 1;5�_�                    )   ,    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�(     �   (   *   ?      -                     if bitCounter = 1 then ;5�_�                    )   +    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�)     �   (   *   ?      ,                     if bitCounter = 1 then 5�_�                    *       ����                                                                                                                                                                                                                                                                                                                                                  V        ^�*     �   )   +          C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);5�_�                    *   %    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�1     �   )   +   ?      F                        m_axis_tdata(bitCounter)   <= s_axis_tdata(0);5�_�                    *   /    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�9     �   )   +   ?      P                        m_axis_tdata(7 downto 0bitCounter)   <= s_axis_tdata(0);5�_�                    *   1    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�;     �   )   +   ?      F                        m_axis_tdata(7 downto 0)   <= s_axis_tdata(0);5�_�                    *   1    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�;     �   )   +   ?      E                        m_axis_tdata(7 downto 0)  <= s_axis_tdata(0);5�_�                    *   @    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�?     �   )   +   ?      D                        m_axis_tdata(7 downto 0) <= s_axis_tdata(0);5�_�                    *   @    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�?     �   )   +   ?      C                        m_axis_tdata(7 downto 0) <= s_axis_tdata0);5�_�                    *   @    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�?     �   )   +   ?      B                        m_axis_tdata(7 downto 0) <= s_axis_tdata);5�_�                    +   *    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�B     �   *   ,   ?    �   +   ,   ?    5�_�                    +       ����                                                                                                                                                                                                                                                                                                                                                  V        ^�D     �   *   ,   @      +                     if bitCounter = 1 then5�_�                    +       ����                                                                                                                                                                                                                                                                                                                                                  V        ^�I     �   *   ,   @    �   +   ,   @    5�_�                    +        ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�J     �   *   ,          B                     bitCounter                 := bitCounter + 1;5�_�                   *        ����                                                                                                                                                                                                                                                                                                                            +           *           V        ^�Q     �   >   @   A         end process shift_reg;�   =   ?   A            end if;�   <   >   A               end if;�   ;   =   A                  end case;�   :   <   A                        end if;�   9   ;   A      7                        state         <= waitingSvalid;�   8   :   A      +                        bitCounter    := 0;�   7   9   A      -                        s_axis_tready <= '1';�   6   8   A      -                        m_axis_tvalid <= '0';�   5   7   A      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   4   6   A      $               when waitingMready =>�   3   5   A                        end if;�   2   4   A                           end if;�   1   3   A      7                        state         <= waitingMready;�   0   2   A      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   /   1   A      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   .   0   A      \                     if bitCounter = 8 then                             --porque bit voy?   �   -   /   A      B                     bitCounter                 := bitCounter + 1;�   ,   .   A      C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);�   +   -   A      3                        elsewif bitCounter = 1 then�   *   ,   A      C                        bitCounter               := bitCounter + 1;�   )   +   A      A                        m_axis_tdata(7 downto 0) <= s_axis_tdata;�   (   *   A      +                     if bitCounter = 1 then�   '   )   A      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   A      $               when waitingSvalid =>�   %   '   A                  case state is�   $   &   A               else�   #   %   A                  bitCounter    := 0;�   "   $   A      -            m_axis_tdata  <= (others => '0');�   !   #   A      !            m_axis_tvalid <= '0';�       "   A      !            s_axis_tready <= '1';�      !   A      +            state         <= waitingSvalid;�          A               if rst = '0' then�         A            if rising_edge(clk) then�         A         begin�         A      0      variable bitCounter :integer range 0 to 8;�         A         shift_reg:process (clk) is�         A      ,   signal state:shiftState := waitingSvalid;�         A      *           rst           : in  STD_LOGIC);�         A      )           clk           : in  STD_LOGIC;�         A      )           s_axis_tready : out STD_LOGIC;�         A      )           s_axis_tlast  : in  STD_LOGIC;�         A      )           s_axis_tvalid : in  STD_LOGIC;�         A      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      A      )           m_axis_tready : in  STD_LOGIC;�   	      A      )           m_axis_tlast  : out STD_LOGIC;�      
   A      )           m_axis_tvalid : out STD_LOGIC;�      	   A      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�         A          Port(  �   )   +          A                        m_axis_tdata(7 downto 0) <= s_axis_tdata;�   *   ,          E                        bitCounter                 := bitCounter + 1;5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                            +           *           V        ^�U     �   +   .   A      3                        elsewif bitCounter = 1 then5�_�                    )   %    ����                                                                                                                                                                                                                                                                                                                            +           *           V        ^�Z     �   (   *   B      +                     if bitCounter = 1 then5�_�                    -        ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^�_     �   ,   /   A    �   -   .   A    �   ,   -          2                           wif bitCounter = 1 then5�_�                     -   %    ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�b     �   ,   .   C      A                        m_axis_tdata(7 downto 0) <= s_axis_tdata;5�_�      !               -   /    ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�h     �   ,   .   C      B                        m_axis_tdata(15 downto 0) <= s_axis_tdata;5�_�       "           !   .   4    ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�r     �   -   /   C      C                        bitCounter               := bitCounter + 1;5�_�   !   #           "   .   4    ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�s     �   -   /   C      4                        bitCounter               := 5�_�   "   $           #   /       ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�w     �   .   /          C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);5�_�   #   %           $   /       ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�x     �   .   /          B                     bitCounter                 := bitCounter + 1;5�_�   $   &           %   /       ����                                                                                                                                                                                                                                                                                                                            -           .   B       V        ^�y     �   .   /          \                     if bitCounter = 8 then                             --porque bit voy?   5�_�   %   '           &   0        ����                                                                                                                                                                                                                                                                                                                            0   "       0   "       V   "    ^�|     �   /   0          `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�   &   (           '   /       ����                                                                                                                                                                                                                                                                                                                            0   "       0   "       V   "    ^�}     �   .   0   ?    �   /   0   ?    5�_�   '   )           (   -        ����                                                                                                                                                                                                                                                                                                                            -   *       1   *       V   *    ^�     �   0   2          7                        state         <= waitingMready;�   /   1          l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   .   0          `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   -   /          6                        bitCounter               := 0;�   ,   .          B                        m_axis_tdata(15 downto 8) <= s_axis_tdata;5�_�   (   *           )   .       ����                                                                                                                                                                                                                                                                                                                            -   *       1   *       V   *    ^�     �   -   .          9                           bitCounter               := 0;5�_�   )   +           *   -        ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�    �   <   >   ?         end process shift_reg;�   ;   =   ?            end if;�   :   <   ?               end if;�   9   ;   ?                  end case;�   8   :   ?                        end if;�   7   9   ?      7                        state         <= waitingSvalid;�   6   8   ?      +                        bitCounter    := 0;�   5   7   ?      -                        s_axis_tready <= '1';�   4   6   ?      -                        m_axis_tvalid <= '0';�   3   5   ?      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   2   4   ?      $               when waitingMready =>�   1   3   ?                        end if;�   0   2   ?                           end if;�   /   1   ?      F                           state                     <= waitingMready;�   .   0   ?      {                           s_axis_tready             <= '0';                              --entonces yo tambien estoy listo�   -   /   ?      o                           m_axis_tvalid             <= '1';                           --y ya no tengo mas nada�   ,   .   ?      E                           m_axis_tdata(15 downto 8) <= s_axis_tdata;�   +   -   ?                              else �   *   ,   ?      C                        bitCounter               := bitCounter + 1;�   )   +   ?      A                        m_axis_tdata(7 downto 0) <= s_axis_tdata;�   (   *   ?      +                     if bitCounter = 0 then�   '   )   ?      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   ?      $               when waitingSvalid =>�   %   '   ?                  case state is�   $   &   ?               else�   #   %   ?                  bitCounter    := 0;�   "   $   ?      -            m_axis_tdata  <= (others => '0');�   !   #   ?      !            m_axis_tvalid <= '0';�       "   ?      !            s_axis_tready <= '1';�      !   ?      +            state         <= waitingSvalid;�          ?               if rst = '0' then�         ?            if rising_edge(clk) then�         ?         begin�         ?      0      variable bitCounter :integer range 0 to 8;�         ?         shift_reg:process (clk) is�         ?      ,   signal state:shiftState := waitingSvalid;�         ?      *           rst           : in  STD_LOGIC);�         ?      )           clk           : in  STD_LOGIC;�         ?      )           s_axis_tready : out STD_LOGIC;�         ?      )           s_axis_tlast  : in  STD_LOGIC;�         ?      )           s_axis_tvalid : in  STD_LOGIC;�         ?      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      ?      )           m_axis_tready : in  STD_LOGIC;�   	      ?      )           m_axis_tlast  : out STD_LOGIC;�      
   ?      )           m_axis_tvalid : out STD_LOGIC;�      	   ?      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�         ?          Port(  �   ,   .          E                           m_axis_tdata(15 downto 8) <= s_axis_tdata;�   /   1          :                           state         <= waitingMready;�   .   0          o                           s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   -   /          c                           m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      W--junto 8 bytes en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   +   -           ,      
    ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      Y--junto 168 bytes en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      X--junto 16 bytes en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      X--junto 16 bites en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      W--junto 16 bits en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�     �         ?      b--junto 2 bytes de 8  bits en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                            -          0          V       ^�    �         ?      --junto 2 bytes de 8  5�_�   1   3           2           ����                                                                                                                                                                                                                                                                                                                                                  V        ^$     �         ?    �         ?    5�_�   2   6           3          ����                                                                                                                                                                                                                                                                                                                                                  V        ^$     �         C    5�_�   3   7   5       6          ����                                                                                                                                                                                                                                                                                                                                                       ^$     �         D      )           m_axis_tvalid : out STD_LOGIC;   )           m_axis_tlast  : out STD_LOGIC;   )           m_axis_tready : in  STD_LOGIC;�         D      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);5�_�   6   8           7      8    ����                                                                                                                                                                                                                                                                                                                                                       ^$     �         D      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (15 downto 0);5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                       ^$      �                0           m_axis_config_tlast  : out STD_LOGIC;5�_�   8   @           9           ����                                                                                                                                                                                                                                                                                                                                      A          V       ^$/     �   @   B   C         end process shift_reg;�          C         shift_reg:process (clk) is5�_�   9   A   :       @   B        ����                                                                                                                                                                                                                                                                                                                                      A          V       ^$k     �   A   E   C    �   B   C   C    5�_�   @   B           A   B        ����                                                                                                                                                                                                                                                                                                                                      A          V       ^$m     �   A   C   F    5�_�   A   C           B   C        ����                                                                                                                                                                                                                                                                                                                            C          D          V       ^$p     �   B   D   G      #m_axis_config_tdata  <= "00000001";�   @   B   G          end process shift_reg;/*}}}*/�   ?   A   G            end if;�   >   @   G               end if;�   =   ?   G                  end case;�   <   >   G                        end if;�   ;   =   G      7                        state         <= waitingSvalid;�   :   <   G      +                        bitCounter    := 0;�   9   ;   G      -                        s_axis_tready <= '1';�   8   :   G      -                        m_axis_tvalid <= '0';�   7   9   G      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   6   8   G      $               when waitingMready =>�   5   7   G                        end if;�   4   6   G                           end if;�   3   5   G      F                           state                     <= waitingMready;�   2   4   G      {                           s_axis_tready             <= '0';                              --entonces yo tambien estoy listo�   1   3   G      o                           m_axis_tvalid             <= '1';                           --y ya no tengo mas nada�   0   2   G      E                           m_axis_tdata(15 downto 8) <= s_axis_tdata;�   /   1   G                              else �   .   0   G      C                        bitCounter               := bitCounter + 1;�   -   /   G      A                        m_axis_tdata(7 downto 0) <= s_axis_tdata;�   ,   .   G      +                     if bitCounter = 0 then�   +   -   G      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   *   ,   G      $               when waitingSvalid =>�   )   +   G                  case state is�   (   *   G               else�   '   )   G                  bitCounter    := 0;�   &   (   G      -            m_axis_tdata  <= (others => '0');�   %   '   G      !            m_axis_tvalid <= '0';�   $   &   G      !            s_axis_tready <= '1';�   #   %   G      +            state         <= waitingSvalid;�   "   $   G               if rst = '0' then�   !   #   G            if rising_edge(clk) then�       "   G         begin�      !   G      0      variable bitCounter :integer range 0 to 8;�          G      $   shift_reg:process (clk) is/*{{{*/�         G      ,   signal state:shiftState := waitingSvalid;�         G      *           rst           : in  STD_LOGIC);�         G      )           clk           : in  STD_LOGIC;�         G      0           m_axis_config_tready : in  STD_LOGIC;�         G      0           m_axis_config_tvalid : out STD_LOGIC;�         G      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (8 downto 0);�         G      )           s_axis_tready : out STD_LOGIC;�         G      )           s_axis_tlast  : in  STD_LOGIC;�         G      )           s_axis_tvalid : in  STD_LOGIC;�         G      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      G      )           m_axis_tready : in  STD_LOGIC;�   	      G      )           m_axis_tlast  : out STD_LOGIC;�      
   G      )           m_axis_tvalid : out STD_LOGIC;�      	   G      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�         G          Port(  �         G       --junto 2 bytes de 8  en 1 de 16�   B   D          #m_axis_config_tdata <= "00000001"; �   C   E          m_axis_config_tvalid <= '1';5�_�   B   D           C   E        ����                                                                                                                                                                                                                                                                                                                            C          D          V       ^$q    �   D   E          m_axis_config_tready 5�_�   C   E           D           ����                                                                                                                                                                                                                                                                                                                                                             ^$�     �   @   B   F          end process shift_reg;/*}}}*/�          F      $   shift_reg:process (clk) is/*{{{*/5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                  V        ^$�     �          F      !   shift_reg:process (clk) is/**/5�_�   E   G           F   A       ����                                                                                                                                                                                                                                                                                                                                                  V        ^$�     �   @   B   F         end process shift_reg;/**/5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$�    �   @   B   F         end process shift_reg;�          F         shift_reg:process (clk) is5�_�   G   I           H      8    ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$�   	 �         F      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (8 downto 0);5�_�   H   J           I   D       ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$"N     �   C   E   F      m_axis_config_tvalid <= '1';5�_�   I   K           J   D   (    ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$"Z   
 �   C   E   F      ,m_axis_config_tvalid <= '1'; --inverse IDFTT5�_�   J   L           K   D       ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$"m     �   C   E   F      +m_axis_config_tvalid <= '1'; --inverse IFTT5�_�   K   M           L   C   "    ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$"n     �   B   D   F      #m_axis_config_tdata  <= "00000001";�   C   D   F    5�_�   L   N           M   C   #    ����                                                                                                                                                                                                                                                                                                                            A                    V       ^$"q    �   B   D   F      1m_axis_config_tdata  <= "00000001";--inverse IFTT5�_�   M               N   C        ����                                                                                                                                                                                                                                                                                                                                                             ^-�'    �   B   D   F      2m_axis_config_tdata  <= "00000001"; --inverse IFTT5�_�   9   ;       @   :   B        ����                                                                                                                                                                                                                                                                                                                                                       ^$1     �   A   C   C           5�_�   :   <           ;   C        ����                                                                                                                                                                                                                                                                                                                                                       ^$;     �   C   D   D    �   B   E          m_axis_config_tdata     $m_axis_config_tvalid end Behavioral;   m_axis_config_tready 5�_�   ;   =           <   D       ����                                                                                                                                                                                                                                                                                                                                                       ^$B     �   C   E   E      m_axis_config_tvalid ;5�_�   <   >           =   D       ����                                                                                                                                                                                                                                                                                                                                                       ^$D     �   C   E   E      m_axis_config_tvalid <= '1';5�_�   =   ?           >   C       ����                                                                                                                                                                                                                                                                                                                            C          E          V       ^$Q     �   B   D   E      #m_axis_config_tdata <= "00000001"; 5�_�   >               ?   E        ����                                                                                                                                                                                                                                                                                                                            C           C           V        ^$]     �   D   F        5�_�   3       4   6   5           ����                                                                                                                                                                                                                                                                                                                                                  V        ^$     �              5�_�   3           5   4           ����                                                                                                                                                                                                                                                                                                                                                  V        ^$     �         D      lkk5�_�                    +        ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�L     �   *   ,   A      Ekkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5��