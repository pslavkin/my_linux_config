Vim�UnDo� 6[ނ8>�z�����p�Z�:nGo���}���   Q                                   ]��f    _�                             ����                                                                                                                                                                                                                                                                                                                                                             ]��E     �         :    �         :    5�_�                    %        ����                                                                                                                                                                                                                                                                                                                                                             ]��S     �   $   0   <    �   %   &   <    5�_�                    G        ����                                                                                                                                                                                                                                                                                                                                                             ]��e    �   F   Q   G    �   G            5�_�                    0        ����                                                                                                                                                                                                                                                                                                                                                             ]��_     �   0   1   G    �   /   0   G   
   aaa: component lab1      generic map (                     N => 4                  )      port map (                  clk=>clk_1,                  rst=>reset_rtl,                  swt=>swt_rtl,                  led=>led_rtl               );5��