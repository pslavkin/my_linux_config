Vim�UnDo� %ỳ�Đ�s��^c�eH�ANT�T����?�H   >   )           n_axis_tready : in  STD_LOGIC;                             ^��    _�                     )        ����                                                                                                                                                                                                                                                                                                                            )          +          V       ^��     �   (   )          C                     --m_axis_tdata(bitCounter) <= s_axis_tdata(0);   B                     --bitCounter               := bitCounter + 1;   B                     --bitCounter               := bitCounter + 1;5�_�                    )        ����                                                                                                                                                                                                                                                                                                                            )          +          V       ^��    �   ;   =   >         end process shift_reg;�   :   <   >            end if;�   9   ;   >               end if;�   8   :   >                  end case;�   7   9   >                        end if;�   6   8   >      7                        state         <= waitingSvalid;�   5   7   >      +                        bitCounter    := 0;�   4   6   >      -                        s_axis_tready <= '1';�   3   5   >      -                        m_axis_tvalid <= '0';�   2   4   >      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   1   3   >      $               when waitingMready =>�   0   2   >                        end if;�   /   1   >                           end if;�   .   0   >      7                        state         <= waitingMready;�   -   /   >      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   ,   .   >      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   +   -   >      \                     if bitCounter = 8 then                             --porque bit voy?   �   *   ,   >      B                     bitCounter                 := bitCounter + 2;�   )   +   >      C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);�   (   *   >      C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);�   '   )   >      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   >      $               when waitingSvalid =>�   %   '   >                  case state is�   $   &   >               else�   #   %   >                  bitCounter    := 0;�   "   $   >      -            m_axis_tdata  <= (others => '0');�   !   #   >      !            m_axis_tvalid <= '0';�       "   >      !            s_axis_tready <= '1';�      !   >      +            state         <= waitingSvalid;�          >               if rst = '0' then�         >            if rising_edge(clk) then�         >         begin�         >      0      variable bitCounter :integer range 0 to 8;�         >         shift_reg:process (clk) is�         >      ,   signal state:shiftState := waitingSvalid;�         >      5   type shiftState is (waitingSvalid, waitingMready);�         >      *           rst           : in  STD_LOGIC);�         >      )           clk           : in  STD_LOGIC;�         >      )           s_axis_tready : out STD_LOGIC;�         >      )           s_axis_tlast  : in  STD_LOGIC;�         >      )           s_axis_tvalid : in  STD_LOGIC;�         >      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      >      )           n_axis_tready : in  STD_LOGIC;�   	      >      )           m_axis_tlast  : out STD_LOGIC;�      
   >      )           m_axis_tvalid : out STD_LOGIC;�      	   >      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         >          Port(  �   (   *          C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);�   *   ,          @                     bitCounter               := bitCounter + 2;�   )   +          C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);5�_�                            ����                                                                                                                                                                                                                                                                                                                            )          +          V       ^��     �         >      5   type shiftState is (waitingSvalid, waitingMready);5�_�                            ����                                                                                                                                                                                                                                                                                                                            )          +          V       ^��    �         >      2type shiftState is (waitingSvalid, waitingMready);5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ^�e    �                'architecture Behavioral of join_8to1 is�                end join_8to1;�                entity join_8to1 is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   
      >      )           n_axis_tready : in  STD_LOGIC;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   
      >      )           m_axis_tready : in  STD_LOGIC;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   
      >      )           n_axis_tready : in  STD_LOGIC;5��