Vim�UnDo� �CWA�|�r)H3������*iS����y*�   L   D                        index         := to_integer(unsigned(test));   2   =     �      �  �  �    ^V�   t _�                             ����                                                                                                                                                                                                                                                                                                                                                v       ^�5     �                'architecture Behavioral of join_8to1 is�                end join_8to1;�                entity join_8to1 is5�_�                    )   !    ����                                                                                                                                                                                                                                                                                                                            )   !       )   ,       v   ,    ^�N     �   (   *   =      A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);5�_�                    )   1    ����                                                                                                                                                                                                                                                                                                                            )   !       )   ,       v   ,    ^�P     �   (   *   =      5                     m_axis_tdata <= s_axis_tdata(0);5�_�                    )   1    ����                                                                                                                                                                                                                                                                                                                            )   !       )   ,       v   ,    ^�P     �   (   *   =      4                     m_axis_tdata <= s_axis_tdata0);5�_�                    )   1    ����                                                                                                                                                                                                                                                                                                                            )   !       )   ,       v   ,    ^�Q     �   (   *   =      3                     m_axis_tdata <= s_axis_tdata);5�_�                    +   %    ����                                                                                                                                                                                                                                                                                                                            )   !       )   ,       v   ,    ^�h     �   *   ,   =      \                     if bitCounter = 8 then                             --porque bit voy?   5�_�      	             )        ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^��     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      7                        state         <= waitingSvalid;�   4   6   =      +                        bitCounter    := 0;�   3   5   =      -                        s_axis_tready <= '1';�   2   4   =      -                        m_axis_tvalid <= '0';�   1   3   =      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   0   2   =      $               when waitingMready =>�   /   1   =                        end if;�   .   0   =                           end if;�   -   /   =      7                        state         <= waitingMready;�   ,   .   =      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   +   -   =      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   *   ,   =      \                     if bitCounter = 1 then                             --porque bit voy?   �   )   +   =      4                     bitCounter   := bitCounter + 1;�   (   *   =      2                     m_axis_tdata <= s_axis_tdata;�   '   )   =      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   =      $               when waitingSvalid =>�   %   '   =                  case state is�   $   &   =               else�   #   %   =                  bitCounter    := 0;�   "   $   =      -            m_axis_tdata  <= (others => '0');�   !   #   =      !            m_axis_tvalid <= '0';�       "   =      !            s_axis_tready <= '1';�      !   =      +            state         <= waitingSvalid;�          =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      =      )           m_axis_tready : in  STD_LOGIC;�   	      =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   (   *          2                     m_axis_tdata <= s_axis_tdata;�   )   +          @                     bitCounter               := bitCounter + 1;5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^�     �         =       5�_�   	              
           ����                                                                                                                                                                                                                                                                                                                            +   %       ,   %       V   %    ^�     �         ?       5�_�   
                    &    ����                                                                                                                                                                                                                                                                                                                            +   %       ,   %       V   %    ^��     �         ?      ,type mapp_table is array (15 to 0) of signed5�_�                       &    ����                                                                                                                                                                                                                                                                                                                            +   %       ,   %       V   %    ^��     �         ?      &type mapp_table is array (15 to 0) of 5�_�                       
    ����                                                                                                                                                                                                                                                                                                                            ,   %       -   %       V   %    ^�-     �         @      ?type mapp_table is array (15 to 0) of integer range -128 to 1275�_�                       ?    ����                                                                                                                                                                                                                                                                                                                            ,   %       -   %       V   %    ^�1     �         @      ?type mapp_array is array (15 to 0) of integer range -128 to 1275�_�                       ?    ����                                                                                                                                                                                                                                                                                                                            ,   %       -   %       V   %    ^�2     �         @    5�_�                           ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^�5     �         A      @type mapp_array is array (15 to 0) of integer range -128 to 127;5�_�                           ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^�7     �         A      ?type map_array is array (15 to 0) of integer range -128 to 127;5�_�                            ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^�J     �         A       5�_�                       #    ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^��     �         A      'signal mapper_table : mapper_array := (5�_�                       '    ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^��    �         A      'signal mapper_table : mapper_array <= (5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^�)    �         A      -signal mapper_table : mapper_array <= (0=>1);5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                            -   %       .   %       V   %    ^�t    �         A      ,signal mapper_table : mapper_array <= (0=>1)5�_�                            ����                                                                                                                                                                                                                                                                                                                               ,          ,       V   ,    ^�     �                -signal mapper_table : mapper_array <= (0=>1);5�_�                            ����                                                                                                                                                                                                                                                                                                                               ,          ,       V   ,    ^�     �         @    �         @    5�_�                            ����                                                                                                                                                                                                                                                                                                                               ,          ,       V   ,    ^�    �                -signal mapper_table : mapper_array <= (0=>1);5�_�                           ����                                                                                                                                                                                                                                                                                                                               ,          ,       V   ,    ^�     �         A      ,   signal state:shiftState := waitingSvalid;5�_�                           ����                                                                                                                                                                                                                                                                                                                               ,          ,       V   ,    ^�    �         A      4   signal state        :shiftState := waitingSvalid;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �                Btype mapper_array is array (15 to 0) of integer range -128 to 127;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         @    �         @    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         B       �         A    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �                   k5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                                V       ^�    �                Btype mapper_array is array (15 to 0) of integer range -128 to 127;5�_�       "           !      &    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         A      0   signal mapper_table : mapper_array <= (0=>1);5�_�   !   #           "      '    ����                                                                                                                                                                                                                                                                                                                                                V       ^�    �         A      1   signal mapper_table : mapper_array :<= (0=>1);5�_�   "   $           #      -    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         A      0   signal mapper_table : mapper_array := (0=>1);5�_�   #   %           $      /    ����                                                                                                                                                                                                                                                                                                                                                V       ^��    �         A      1   signal mapper_table : mapper_array := (0=>"1);5�_�   $   &           %      -    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      2   signal mapper_table : mapper_array := (0=>"1");5�_�   %   '           &      .    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      1   signal mapper_table : mapper_array := (0=>1");5�_�   &   (           '      -    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      0   signal mapper_table : mapper_array := (0=>1);5�_�   '   )           (      0    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      3   signal mapper_table : mapper_array := (0=>1231);5�_�   (   *           )      -    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      2   signal mapper_table : mapper_array := (0=>123);5�_�   )   +           *      1    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         A      4   signal mapper_table : mapper_array := (0=>x"123);5�_�   *   -           +      1    ����                                                                                                                                                                                                                                                                                                                                                V       ^��   	 �         A      3   signal mapper_table : mapper_array := (0=>x"12);5�_�   +   .   ,       -      )    ����                                                                                                                                                                                                                                                                                                                                                V       ^�9     �         A      4   signal mapper_table : mapper_array := (0=>x"12");5�_�   -   /           .      4    ����                                                                                                                                                                                                                                                                                                                                                V       ^�A     �         A      ?   signal mapper_table : mapper_array := "1","2","3"(0=>x"12");5�_�   .   0           /      4    ����                                                                                                                                                                                                                                                                                                                                                V       ^�B   
 �         A      4   signal mapper_table : mapper_array := "1","2","3"5�_�   /   1           0      ,    ����                                                                                                                                                                                                                                                                                                                                                V       ^�L    �         A      5   signal mapper_table : mapper_array := "1","2","3";5�_�   0   2           1      )    ����                                                                                                                                                                                                                                                                                                                                                V       ^�[     �         A      -   signal mapper_table : mapper_array := "1";5�_�   1   3           2      *    ����                                                                                                                                                                                                                                                                                                                                                V       ^�\    �         A      ,   signal mapper_table : mapper_array := 1";5�_�   2   4           3      *    ����                                                                                                                                                                                                                                                                                                                                                V       ^�e    �         A      +   signal mapper_table : mapper_array := 1;5�_�   3   5           4      )    ����                                                                                                                                                                                                                                                                                                                                                V       ^�y     �         A      P   signal mapper_table : mapper_array := 1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16;5�_�   4   6           5      P    ����                                                                                                                                                                                                                                                                                                                                                V       ^�|    �         A      Q   signal mapper_table : mapper_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16;5�_�   5   7           6      M    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         A      R   signal mapper_table : mapper_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16);5�_�   6   8           7      M    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         A      Q   signal mapper_table : mapper_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,1516);5�_�   7   9           8      M    ����                                                                                                                                                                                                                                                                                                                                                V       ^�    �         A      P   signal mapper_table : mapper_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,156);5�_�   8   :           9      2    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�    �         A      E   type mapper_array is array (15 to 0) of integer range -128 to 127;5�_�   9   ;           :      )    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^��     �         A      O   signal mapper_table : mapper_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,15);5�_�   :   <           ;      )    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^��    �         A      )   signal mapper_table : mapper_array := 5�_�   ;   =           <      *    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^��    �         A      7   signal mapper_table : mapper_array := (others => 0);5�_�   <   >           =      *    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         A      ;   signal mapper_table : mapper_array := (1,2,others => 0);5�_�   =   ?           >      /    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�    �         A      >   signal mapper_table : mapper_array := (0=>1,2,others => 0);5�_�   >   @           ?      +    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         A      A   signal mapper_table : mapper_array := (0=>1,1=>2,others => 0);5�_�   ?   A           @      ,    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         A      C   signal mapper_table : mapper_array := (0 l=>1,1=>2,others => 0);5�_�   @   B           A      .    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         A      B   signal mapper_table : mapper_array := (0 =>1,1=>2,others => 0);5�_�   A   C           B      2    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         A      C   signal mapper_table : mapper_array := (0 => 1,1=>2,others => 0);5�_�   B   D           C      5    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�    �         A      D   signal mapper_table : mapper_array := (0 => 1,1 =>2,others => 0);5�_�   C   E           D      /    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�      �         A    5�_�   D   F           E      /    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�$     �         B      E   signal mapper_table : mapper_array := (0 => 1,1 => 2,others => 0);5�_�   E   G           F      1    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�%     �         B      F   signal mapper_table : mapper_array := (0 => "1,1 => 2,others => 0);5�_�   F   H           G      8    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�'     �         B      G   signal mapper_table : mapper_array := (0 => "1",1 => 2,others => 0);5�_�   G   I           H      :    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�)    �         B      H   signal mapper_table : mapper_array := (0 => "1",1 => "2,others => 0);5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^��     �         B      I   signal mapper_table : mapper_array := (0 => "1",1 => "2",others => 0);5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^��     �         B      L   constant  mapper_table : mapper_array := (0 => "1",1 => "2",others => 0);5�_�   J   L           K      1    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         B      K   constant mapper_table : mapper_array := (0 => "1",1 => "2",others => 0);5�_�   K   M           L      2    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         B      J   constant mapper_table : mapper_array := (0 => 1",1 => "2",others => 0);5�_�   L   N           M      8    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�     �         B      I   constant mapper_table : mapper_array := (0 => 1,1 => "2",others => 0);5�_�   M   O           N      9    ����                                                                                                                                                                                                                                                                                                                               2          C       v   C    ^�    �         B      H   constant mapper_table : mapper_array := (0 => 1,1 => 2",others => 0);5�_�   N   P           O      ,    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�    �         B      G   constant mapper_table : mapper_array := (0 => 1,1 => 2,others => 0);5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�1     �         B      3   type mapper_array is array (15 to 0) of integer;5�_�   P   R           Q      $    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�4     �         B      2   type mapper_array is array (0 to 0) of integer;5�_�   Q   S           R      &    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�5    �         B      4   type mapper_array is array (0 to 150) of integer;5�_�   R   T           S      ,    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�:    �         B      9   constant mapper_table : mapper_array := (others => 0);5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�]     �         B      3   type mapper_array is array (0 to 15) of integer;5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         B    �         B    5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         C      1   type real_array is array (0 to 15) of integer;5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         C      /   type im_array is array (0 to 15) of integer;5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         C      =   constant mapper_table : mapper_array := (1,2,others => 0);5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         C      ;   constant real_table : mapper_array := (1,2,others => 0);5�_�   Y   [           Z      '    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �          C      9   constant real_table : real_array := (1,2,others => 0);5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �      .   E         �         E    5�_�   [   ]           \           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         T         1255�_�   \   ^           ]           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         T        1255�_�   ]   _           ^           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         T       1255�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         T      1255�_�   _   a           `          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         T      125,   1065�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         S      	125, 106,   71�         S      125, 1065�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         R      125, 106, 71,   25�         R      125, 106, 715�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         Q      125, 106, 71, 25,   -25�         Q      125, 106, 71, 255�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         P      125, 106, 71, 25, -25,   -71�         P      125, 106, 71, 25, -255�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         O      125, 106, 71, 25, -25, -71,   -106�         O      125, 106, 71, 25, -25, -715�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         N      !125, 106, 71, 25, -25, -71, -106,   -125�         N       125, 106, 71, 25, -25, -71, -1065�_�   f   h           g      &    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         M      '125, 106, 71, 25, -25, -71, -106, -125,   -125�         M      &125, 106, 71, 25, -25, -71, -106, -1255�_�   g   i           h      ,    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         L      -125, 106, 71, 25, -25, -71, -106, -125, -125,   -106�         L      ,125, 106, 71, 25, -25, -71, -106, -125, -1255�_�   h   j           i      2    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         K      3125, 106, 71, 25, -25, -71, -106, -125, -125, -106,   -71�         K      2125, 106, 71, 25, -25, -71, -106, -125, -125, -1065�_�   i   k           j      7    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         J      8125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71,   -25�         J      7125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -715�_�   j   l           k      <    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         I      =125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25,   25�         I      <125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -255�_�   k   m           l      @    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         H      A125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25,   71�         H      @125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 255�_�   l   n           m      D    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^��     �         G      E125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71,   106�         G      D125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 715�_�   m   o           n      I    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�      �         F      J125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106,   125�         F      I125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 1065�_�   n   p           o      N    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         E      N125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 1255�_�   o   q           p      &    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         E      '   constant real_table : real_array :=    P125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   p   r           q      '    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         D      w   constant real_table : real_array := 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�	     �                   (1,2,others => 0);5�_�   r   t           s           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         C    �         C    5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         D      x   constant real_table : real_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         D      v   constant im_table : real_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         D      t   constant im_table : im_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   v   x           w      %    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�     �         D      v   constant im_table   : im_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);5�_�   w   y           x      $    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�      �          D    5�_�   x   z           y           ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�!     �      /   E       �          E    5�_�   y   {           z          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�#     �          T      25,   71�          T      255�_�   z   |           {          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�#     �          S      25, 71,   106�          S      25, 715�_�   {   }           |          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�#     �          R      25, 71, 106,   125�          R      25, 71, 1065�_�   |   ~           }          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          Q      25, 71, 106, 125,   125�          Q      25, 71, 106, 1255�_�   }              ~          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          P      25, 71, 106, 125, 125,   106�          P      25, 71, 106, 125, 1255�_�   ~   �                     ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          O      25, 71, 106, 125, 125, 106,   71�          O      25, 71, 106, 125, 125, 1065�_�      �           �          ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          N      25, 71, 106, 125, 125, 106, 71,   25�          N      25, 71, 106, 125, 125, 106, 715�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          M      #25, 71, 106, 125, 125, 106, 71, 25,   -25�          M      "25, 71, 106, 125, 125, 106, 71, 255�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          L      (25, 71, 106, 125, 125, 106, 71, 25, -25,   -71�          L      '25, 71, 106, 125, 125, 106, 71, 25, -255�_�   �   �           �      ,    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          K      -25, 71, 106, 125, 125, 106, 71, 25, -25, -71,   -106�          K      ,25, 71, 106, 125, 125, 106, 71, 25, -25, -715�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          J      325, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106,   -125�          J      225, 71, 106, 125, 125, 106, 71, 25, -25, -71, -1065�_�   �   �           �      8    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          I      925, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125,   -125�          I      825, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -1255�_�   �   �           �      >    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�$     �          H      ?25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125,   -106�          H      >25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -1255�_�   �   �           �      D    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�%     �          G      E25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106,   -71�          G      D25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -1065�_�   �   �           �      I    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�%     �          F      J25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71,   -25�          F      I25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -715�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�'     �         E      %   constant im_table   : im_array :=    N25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -255�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�(     �         D      s   constant im_table   : im_array := 25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -255�_�   �   �           �      t    ����                                                                                                                                                                                                                                                                                                                               ,          9       v   9    ^�+     �         D      t   constant im_table   : im_array := (25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -255�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               u          u       V   u    ^�/     �   A   C   D         end process shift_reg;�   @   B   D            end if;�   ?   A   D               end if;�   >   @   D                  end case;�   =   ?   D                        end if;�   <   >   D      7                        state         <= waitingSvalid;�   ;   =   D      +                        bitCounter    := 0;�   :   <   D      -                        s_axis_tready <= '1';�   9   ;   D      -                        m_axis_tvalid <= '0';�   8   :   D      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   7   9   D      $               when waitingMready =>�   6   8   D                        end if;�   5   7   D                           end if;�   4   6   D      7                        state         <= waitingMready;�   3   5   D      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   2   4   D      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   1   3   D      \                     if bitCounter = 1 then                             --porque bit voy?   �   0   2   D      4                     bitCounter   := bitCounter + 1;�   /   1   D      2                     m_axis_tdata <= s_axis_tdata;�   .   0   D      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   -   /   D      $               when waitingSvalid =>�   ,   .   D                  case state is�   +   -   D               else�   *   ,   D                  bitCounter    := 0;�   )   +   D      -            m_axis_tdata  <= (others => '0');�   (   *   D      !            m_axis_tvalid <= '0';�   '   )   D      !            s_axis_tready <= '1';�   &   (   D      +            state         <= waitingSvalid;�   %   '   D               if rst = '0' then�   $   &   D            if rising_edge(clk) then�   #   %   D         begin�   "   $   D      0      variable bitCounter :integer range 0 to 8;�   !   #   D         shift_reg:process (clk) is�         D      x   constant im_table   : im_array   := (25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25);�         D      x   constant real_table : real_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);�         D      5   signal state        : shiftState := waitingSvalid;�         D      1   type im_array   is array (0 to 15) of integer;�         D      1   type real_array is array (0 to 15) of integer;�         D      5   type shiftState is (waitingSvalid, waitingMready);�         D      *           rst           : in  STD_LOGIC);�         D      )           clk           : in  STD_LOGIC;�         D      )           s_axis_tready : out STD_LOGIC;�         D      )           s_axis_tlast  : in  STD_LOGIC;�         D      )           s_axis_tvalid : in  STD_LOGIC;�         D      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      D      )           m_axis_tready : in  STD_LOGIC;�   	      D      )           m_axis_tlast  : out STD_LOGIC;�      
   D      )           m_axis_tvalid : out STD_LOGIC;�      	   D      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         D          Port(  �                x   constant real_table : real_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);�                v   constant im_table   : im_array := (25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^�3     �   A   C   D         end process shift_reg;�   @   B   D            end if;�   ?   A   D               end if;�   >   @   D                  end case;�   =   ?   D                        end if;�   <   >   D      7                        state         <= waitingSvalid;�   ;   =   D      +                        bitCounter    := 0;�   :   <   D      -                        s_axis_tready <= '1';�   9   ;   D      -                        m_axis_tvalid <= '0';�   8   :   D      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   7   9   D      $               when waitingMready =>�   6   8   D                        end if;�   5   7   D                           end if;�   4   6   D      7                        state         <= waitingMready;�   3   5   D      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   2   4   D      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   1   3   D      \                     if bitCounter = 1 then                             --porque bit voy?   �   0   2   D      4                     bitCounter   := bitCounter + 1;�   /   1   D      2                     m_axis_tdata <= s_axis_tdata;�   .   0   D      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   -   /   D      $               when waitingSvalid =>�   ,   .   D                  case state is�   +   -   D               else�   *   ,   D                  bitCounter    := 0;�   )   +   D      -            m_axis_tdata  <= (others => '0');�   (   *   D      !            m_axis_tvalid <= '0';�   '   )   D      !            s_axis_tready <= '1';�   &   (   D      +            state         <= waitingSvalid;�   %   '   D               if rst = '0' then�   $   &   D            if rising_edge(clk) then�   #   %   D         begin�   "   $   D      0      variable bitCounter :integer range 0 to 8;�   !   #   D         shift_reg:process (clk) is�         D      �   constant im_table   : im_array   := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         D      �   constant real_table : real_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         D      5   signal state        : shiftState := waitingSvalid;�         D      1   type im_array   is array (0 to 15) of integer;�         D      1   type real_array is array (0 to 15) of integer;�         D      5   type shiftState is (waitingSvalid, waitingMready);�         D      *           rst           : in  STD_LOGIC);�         D      )           clk           : in  STD_LOGIC;�         D      )           s_axis_tready : out STD_LOGIC;�         D      )           s_axis_tlast  : in  STD_LOGIC;�         D      )           s_axis_tvalid : in  STD_LOGIC;�         D      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      D      )           m_axis_tready : in  STD_LOGIC;�   	      D      )           m_axis_tlast  : out STD_LOGIC;�      
   D      )           m_axis_tvalid : out STD_LOGIC;�      	   D      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         D          Port(  �                x   constant real_table : real_array := (125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25, 25, 71, 106, 125);�                x   constant im_table   : im_array   := (25, 71, 106, 125, 125, 106, 71, 25, -25, -71, -106, -125, -125, -106, -71, -25);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^�>     �                5   signal state        : shiftState := waitingSvalid;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^�>    �         C    �         C    5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                               0          0          0    ^�N    �         D      1   type im_array   is array (0 to 15) of integer;�         D      1   type real_array is array (0 to 15) of integer;5�_�   �   �           �      7    ����                                                                                                                                                                                                                                                                                                                               7          7          7    ^�i     �         D      E   type real_array is array (0 to 15) of integer range (-128 to 127);   E   type im_array   is array (0 to 15) of integer range (-128 to 127);5�_�   �   �           �      B    ����                                                                                                                                                                                                                                                                                                                               B          B          B    ^�k    �         D      D   type real_array is array (0 to 15) of integer range -128 to 127);   D   type im_array   is array (0 to 15) of integer range -128 to 127);5�_�   �   �           �   0   1    ����                                                                                                                                                                                                                                                                                                                               B          B          B    ^��     �   0   2   E                           �   0   2   D    5�_�   �   �   �       �   /       ����                                                                                                                                                                                                                                                                                                                               B          B          B    ^��     �   /   1   F                           �   /   1   E    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                               B          B          B    ^��     �   /   1   F      !                     s_axis_tdata5�_�   �   �           �   0        ����                                                                                                                                                                                                                                                                                                                            0           0   +       v   +    ^��     �   /   1   F      8                     real_table(to_unsigned(s_axis_tdata5�_�   �   �           �   0   ,    ����                                                                                                                                                                                                                                                                                                                            0           0   +       v   +    ^��     �   /   1   F      ,                     real_table(s_axis_tdata5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            0          0   -       v   -    ^��     �   /   1   F      .                     real_table(s_axis_tdata);5�_�   �   �           �   1   %    ����                                                                                                                                                                                                                                                                                                                            1   %       1   0       v   0    ^��     �   0   2   F      2                     m_axis_tdata <= s_axis_tdata;�   1   2   F    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            1   %       1   =       v   0    ^��     �   /   0                               5�_�   �   �           �   0   >    ����                                                                                                                                                                                                                                                                                                                            0   %       0   =       v   0    ^��    �   /   1   E      ?                     m_axis_tdata <= real_table(s_axis_tdata);;5�_�   �   �           �   0   0    ����                                                                                                                                                                                                                                                                                                                            0   %       0   =       v   0    ^��     �   /   1   E      >                     m_axis_tdata <= real_table(s_axis_tdata);5�_�   �   �           �   0   H    ����                                                                                                                                                                                                                                                                                                                            0   %       0   =       v   0    ^�    �   /   1   E      J                     m_axis_tdata <= real_table(to_unsigned(s_axis_tdata);5�_�   �   �           �   0   H    ����                                                                                                                                                                                                                                                                                                                            0   %       0   =       v   0    ^�5     �   /   1   E      K                     m_axis_tdata <= real_table(to_unsigned(s_axis_tdata));5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            0   %       0   =       v   0    ^�@     �         E    �         E    5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                            1   %       1   =       v   0    ^�W     �         F      use IEEE.STD_LOGIC_1164.ALL;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ^�]   ! �         F      $use IEEE.numeric_STD_LOGIC_1164.ALL;5�_�   �   �   �       �   1   0    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      M                     m_axis_tdata <= real_table(to_unsigned(s_axis_tdata,4));5�_�   �   �           �   1   0    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      L                     m_axis_tdata <= real_table(o_unsigned(s_axis_tdata,4));5�_�   �   �           �   1   0    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      K                     m_axis_tdata <= real_table(_unsigned(s_axis_tdata,4));5�_�   �   �           �   1   E    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      J                     m_axis_tdata <= real_table(unsigned(s_axis_tdata,4));5�_�   �   �           �   1   E    ����                                                                                                                                                                                                                                                                                                                                                v       ^��   $ �   0   2   F      I                     m_axis_tdata <= real_table(unsigned(s_axis_tdata4));5�_�   �   �   �       �   1   0    ����                                                                                                                                                                                                                                                                                                                                                v       ^�X     �   0   2   F      H                     m_axis_tdata <= real_table(unsigned(s_axis_tdata));5�_�   �   �           �   1   Q    ����                                                                                                                                                                                                                                                                                                                                                v       ^�]   % �   0   2   F      S                     m_axis_tdata <= real_table(to_integer(unsigned(s_axis_tdata));5�_�   �   �           �   1   0    ����                                                                                                                                                                                                                                                                                                                                                v       ^�y   & �   0   2   F      T                     m_axis_tdata <= real_table(to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   3    ����                                                                                                                                                                                                                                                                                                                                                v       ^�~   ' �   0   2   F      Y                     m_axis_tdata <= real_table(1);--to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   %    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      Z                     m_axis_tdata <= real_table(1); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   %    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      \                     m_axis_tdata <= toreal_table(1); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      m                     m_axis_tdata <= STD_LOGIC_VECTOR(toreal_table(1); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      l                     m_axis_tdata <= STD_LOGIC_VECTOR(oreal_table(1); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   C    ����                                                                                                                                                                                                                                                                                                                                                v       ^��   ( �   0   2   F      k                     m_axis_tdata <= STD_LOGIC_VECTOR(real_table(1); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   0   2   F      l                     m_axis_tdata <= STD_LOGIC_VECTOR(real_table(1)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   J    ����                                                                                                                                                                                                                                                                                                                                                v       ^��   ) �   0   2   F      s                     m_axis_tdata <= STD_LOGIC_VECTOR(signed(real_table(1)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                               )          /          /    ^��     �         F      <   type real_array is array (0 to 15) of  range -128 to 127;�         F      C   type real_array is array (0 to 15) of integer range -128 to 127;   C   type im_array   is array (0 to 15) of integer range -128 to 127;5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                            1   6       1   <       v   <    ^��     �   0   2   F      t                     m_axis_tdata <= STD_LOGIC_VECTOR(signed(real_table(1))); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   D    ����                                                                                                                                                                                                                                                                                                                            1   6       1   <       v   <    ^�!   , �   0   2   F      m                     m_axis_tdata <= STD_LOGIC_VECTOR(real_table(1))); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �      )    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�?     �         F      <   type real_array is array (0 to 15) of  range -128 to 127;�         F      B   type real_array is array (0 to 15) of signed range -128 to 127;   B   type im_array   is array (0 to 15) of signed range -128 to 127;5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�E     �   0   2   F      l                     m_axis_tdata <= STD_LOGIC_VECTOR(real_table(1)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   <    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�J     �   0   2   F      t                     m_axis_tdata <= STD_LOGIC_VECTOR(signedd(real_table(1)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   J    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�K   - �   0   2   F      s                     m_axis_tdata <= STD_LOGIC_VECTOR(signed(real_table(1)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   6    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�]     �   0   2   F      t                     m_axis_tdata <= STD_LOGIC_VECTOR(signed(real_table(1))); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   M    ����                                                                                                                                                                                                                                                                                                                               )          .          .    ^�i   . �   0   2   F      w                     m_axis_tdata <= STD_LOGIC_VECTOR(to_signed(real_table(1))); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �   �       �   1   %    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��   / �   0   2   F      y                     m_axis_tdata <= STD_LOGIC_VECTOR(to_signed(real_table(1),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   K    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��     �   0   2   F      y                     m_axis_tdata <= std_logic_vector(to_signed(real_table(1),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   W    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��     �   0   2   F      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(s_axis_tdata1),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   K    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��     �   0   2   F      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(s_axis_tdata),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   K    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��     �   0   2   F      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(unsigned(s_axis_tdata),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   l    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��     �   0   2   F      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(to_integer(unsigned(s_axis_tdata),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   1   m    ����                                                                                                                                                                                                                                                                                                                            1   4       1   %       v   %    ^��   0 �   0   2   F      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(to_integer(unsigned(s_axis_tdata))),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   0   K    ����                                                                                                                                                                                                                                                                                                                            1   K       1   o       v   o    ^�     �   0   2   G                           �   0   2   F    5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            2   K       2   o       v   o    ^�     �   0   2   G                           index := �   1   2   G    5�_�   �   �           �   1   C    ����                                                                                                                                                                                                                                                                                                                            2   K       2   o       v   o    ^�     �   0   2   G      C                     index := to_integer(unsigned(s_axis_tdata)),4)5�_�   �   �           �   $   /    ����                                                                                                                                                                                                                                                                                                                            2   K       2   o       v   o    ^�     �   #   %   G    �   $   %   G    5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            3   K       3   o       v   o    ^�     �   $   &   H      0      variable bitCounter :integer range 0 to 8;5�_�   �   �           �   %   )    ����                                                                                                                                                                                                                                                                                                                            3   K       3   o       v   o    ^�     �   $   &   H      +      variable index :integer range 0 to 8;5�_�   �   �           �   %   +    ����                                                                                                                                                                                                                                                                                                                            3   K       3   o       v   o    ^�     �   $   &   H      -      variable index :integer range 0 to 158;5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            3   K       3   o       v   o    ^�#     �   ,   .   H    �   -   .   H    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            4   K       4   o       v   o    ^�$     �   -   /   I                  bitCounter    := 0;5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            4   K       4   o       v   o    ^�&     �   -   .                      inde    := 0;5�_�   �   �           �   3   K    ����                                                                                                                                                                                                                                                                                                                            3   K       3   n       v   n    ^�7     �   2   4   H      �                     m_axis_tdata <= std_logic_vector(to_signed(real_table(to_integer(unsigned(s_axis_tdata)),4),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   2   5    ����                                                                                                                                                                                                                                                                                                                            3   K       3   n       v   n    ^�<     �   1   3   H    �   2   3   H    5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�=     �   2   4   I      D                     index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�?     �   2   4   I                           index := 5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�C     �   1   3   I      D                     index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�G   1 �   1   3   I      F                     ==index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�L     �   1   3   I      F                     --index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�L     �   1   3   I      E                     -index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�M   2 �   2   4   I                            index := 2;5�_�   �   �           �   2   ?    ����                                                                                                                                                                                                                                                                                                                            4   K       4   n       v   n    ^�_   3 �   1   3   I      D                     index := to_integer(unsigned(s_axis_tdata)),4);5�_�   �   �   �       �   2   ?    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^��     �   1   3   I      C                     index := to_integer(unsigned(s_axis_tdata),4);5�_�   �   �           �   2   ?    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^��   5 �   1   3   I      B                     index := to_integer(unsigned(s_axis_tdata)4);5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^��     �   2   3          "                     --index := 2;5�_�   �   �           �   %   +    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^��     �   $   &   H    �   %   &   H    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      ,      variable index :integer range 0 to 15;5�_�   �   �           �   &   #    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      +      variable real :integer range 0 to 15;5�_�   �   �           �   &   (    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      0      variable real :integer range -128 0 to 15;5�_�   �   �           �   &   (    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      /      variable real :integer range -128  to 15;5�_�   �   �           �   &   ,    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      .      variable real :integer range -128 to 15;5�_�   �   �           �   &   .    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I      0      variable real :integer range -128 to 1275;5�_�   �   �           �   &   .    ����                                                                                                                                                                                                                                                                                                                            3          3   (       v   (    ^��     �   %   '   I    �   &   '   I    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            4          4   (       v   (    ^��     �   %   '   J      /      variable real :integer range -128 to 127;5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            4          4   (       v   (    ^��     �   &   (   J      /      variable real :integer range -128 to 127;5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            4          4   (       v   (    ^��     �   &   (   J      2      variable im_part :integer range -128 to 127;5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            4          4   (       v   (    ^��     �   4   6   J    �   5   6   J    5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            4          4   (       v   (    ^��     �   4   6   K    �   5   6   K    5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            5          5           v        ^��     �   4   6   L      }                     m_axis_tdata <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            5          5           v        ^��     �   4   6   L      q                      <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            5          5           v        ^��     �   4   6   L      q                     e<= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            5          5           v        ^��     �   4   6   L      z                     real_parte<= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            5          5           v        ^��     �   4   6   L      y                     real_part<= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �   �       �   &       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^��     �   %   '   L            variable real_part :;�   %   (   L      4      variable real_part :integer range -128 to 127;   4      variable im_part   :integer range -128 to 127;5�_�   �   �           �   5   Q    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�     �   4   6   L    �   5   6   L    5�_�   �   �           �   6   S    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�     �   5   7   M      z                     real_part <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   5   S    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�     �   4   6   M      z                     real_part <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�     �   5   7   M      S                     real_part <= std_logic_vector(to_signed(real_table(index),8));5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�     �   5   7   M      Q                     im_part <= std_logic_vector(to_signed(real_table(index),8));5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�!     �   4   6   M      S                     real_part <= std_logic_vector(to_signed(real_table(index),8));5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�"     �   5   7   M      Q                     im_part := std_logic_vector(to_signed(real_table(index),8));5�_�   �   �           �   6   =    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�'     �   5   7   M      S                     im_part   := std_logic_vector(to_signed(real_table(index),8));5�_�   �   �           �   7   %    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�/     �   6   8   M      }                     m_axis_tdata <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �              �   7   .    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�5     �   6   8   M      �                     m_axis_tdata <= real_partstd_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �                7   .    ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�6     �   6   8   M      .                     m_axis_tdata <= real_part5�_�                  8       ����                                                                                                                                                                                                                                                                                                                            &          '   2          2    ^�8   6 �   7   8          }                     m_axis_tdata <= std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�                 &   ,    ����                                                                                                                                                                                                                                                                                                                            &   ,       '   ,          ,    ^�P     �   %   (   L      8      variable real_part :std_logic_vector (8 downto 0);   8      variable im_part   :std_logic_vector (8 downto 0);5�_�                 &   ,    ����                                                                                                                                                                                                                                                                                                                            &   ,       '   ,          ,    ^�T   7 �   %   (   L      8      variable real_part :std_logic_vector (8 downto 0);   8      variable im_part   :std_logic_vector (8 downto 0);5�_�                 4   >    ����                                                                                                                                                                                                                                                                                                                            &   ,       '   ,          ,    ^��   8 �   3   5   L      A                     index := to_integer(unsigned(s_axis_tdata));5�_�                 4        ����                                                                                                                                                                                                                                                                                                                            4   I       6   I       V   I    ^��     �   I   K   L         end process shift_reg;�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L                        end if;�   D   F   L      7                        state         <= waitingSvalid;�   C   E   L      +                        bitCounter    := 0;�   B   D   L      -                        s_axis_tready <= '1';�   A   C   L      -                        m_axis_tvalid <= '0';�   @   B   L      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   L      $               when waitingMready =>�   >   @   L                        end if;�   =   ?   L                           end if;�   <   >   L      7                        state         <= waitingMready;�   ;   =   L      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   L      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   L      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   L      4                     bitCounter   := bitCounter + 1;�   7   9   L                           �   6   8   L      /                     m_axis_tdata <= real_part;�   5   7   L      Q                     im_part   := std_logic_vector(to_signed(im_table(index),8));�   4   6   L      S                     real_part := std_logic_vector(to_signed(real_table(index),8));�   3   5   L      Q                     index     := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   L      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   L      $               when waitingSvalid =>�   0   2   L                  case state is�   /   1   L               else�   .   0   L                  bitCounter    := 0;�   -   /   L      -            m_axis_tdata  <= (others => '0');�   ,   .   L      !            m_axis_tvalid <= '0';�   +   -   L      !            s_axis_tready <= '1';�   *   ,   L      +            state         <= waitingSvalid;�   )   +   L               if rst = '0' then�   (   *   L            if rising_edge(clk) then�   '   )   L         begin�   &   (   L      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   L      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   L      ,      variable index :integer range 0 to 15;�   #   %   L      0      variable bitCounter :integer range 0 to 8;�   "   $   L         shift_reg:process (clk) is�          L      5   signal state        : shiftState := waitingSvalid;�         L      �   constant im_table   : im_array   := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         L      �   constant real_table : real_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         L      C   type im_array   is array (0 to 15) of integer range -128 to 127;�         L      C   type real_array is array (0 to 15) of integer range -128 to 127;�         L      5   type shiftState is (waitingSvalid, waitingMready);�         L      *           rst           : in  STD_LOGIC);�         L      )           clk           : in  STD_LOGIC;�         L      )           s_axis_tready : out STD_LOGIC;�         L      )           s_axis_tlast  : in  STD_LOGIC;�         L      )           s_axis_tvalid : in  STD_LOGIC;�         L      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         L      )           m_axis_tready : in  STD_LOGIC;�   
      L      )           m_axis_tlast  : out STD_LOGIC;�   	      L      )           m_axis_tvalid : out STD_LOGIC;�      
   L      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   L          Port(  �   3   5          M                     index := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   5   7          Q                     im_part   := std_logic_vector(to_signed(im_table(index),8));�   4   6          S                     real_part := std_logic_vector(to_signed(real_table(index),8));5�_�                 4        ����                                                                                                                                                                                                                                                                                                                            4           7           V        ^��     �   I   K   L         end process shift_reg;�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L                        end if;�   D   F   L      7                        state         <= waitingSvalid;�   C   E   L      +                        bitCounter    := 0;�   B   D   L      -                        s_axis_tready <= '1';�   A   C   L      -                        m_axis_tvalid <= '0';�   @   B   L      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   L      $               when waitingMready =>�   >   @   L                        end if;�   =   ?   L                           end if;�   <   >   L      7                        state         <= waitingMready;�   ;   =   L      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   L      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   L      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   L      4                     bitCounter   := bitCounter + 1;�   7   9   L                           �   6   8   L      /                     m_axis_tdata <= real_part;�   5   7   L      T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   4   6   L      V                     real_part    := std_logic_vector(to_signed(real_table(index),8));�   3   5   L      T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   L      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   L      $               when waitingSvalid =>�   0   2   L                  case state is�   /   1   L               else�   .   0   L                  bitCounter    := 0;�   -   /   L      -            m_axis_tdata  <= (others => '0');�   ,   .   L      !            m_axis_tvalid <= '0';�   +   -   L      !            s_axis_tready <= '1';�   *   ,   L      +            state         <= waitingSvalid;�   )   +   L               if rst = '0' then�   (   *   L            if rising_edge(clk) then�   '   )   L         begin�   &   (   L      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   L      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   L      ,      variable index :integer range 0 to 15;�   #   %   L      0      variable bitCounter :integer range 0 to 8;�   "   $   L         shift_reg:process (clk) is�          L      5   signal state        : shiftState := waitingSvalid;�         L      �   constant im_table   : im_array   := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         L      �   constant real_table : real_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         L      C   type im_array   is array (0 to 15) of integer range -128 to 127;�         L      C   type real_array is array (0 to 15) of integer range -128 to 127;�         L      5   type shiftState is (waitingSvalid, waitingMready);�         L      *           rst           : in  STD_LOGIC);�         L      )           clk           : in  STD_LOGIC;�         L      )           s_axis_tready : out STD_LOGIC;�         L      )           s_axis_tlast  : in  STD_LOGIC;�         L      )           s_axis_tvalid : in  STD_LOGIC;�         L      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         L      )           m_axis_tready : in  STD_LOGIC;�   
      L      )           m_axis_tlast  : out STD_LOGIC;�   	      L      )           m_axis_tvalid : out STD_LOGIC;�      
   L      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   L          Port(  �   3   5          Q                     index     := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   6   8          /                     m_axis_tdata <= real_part;�   5   7          Q                     im_part   := std_logic_vector(to_signed(im_table(index),8));�   4   6          S                     real_part := std_logic_vector(to_signed(real_table(index),8));5�_�                 K        ����                                                                                                                                                                                                                                                                                                                            4           7           V        ^��     �   J   m   L    �   K   L   L    5�_�    	             K       ����                                                                                                                                                                                                                                                                                                                            4           7           V        ^��     �   J   L   n    5�_�    
          	   L       ����                                                                                                                                                                                                                                                                                                                            4           7           V        ^��     �   K   M   o         shift_reg:process (clk) is5�_�  	            
   L   	    ����                                                                                                                                                                                                                                                                                                                            4           7           V        ^��     �   K   M   o         mapper:process (clk) is5�_�  
               N        ����                                                                                                                                                                                                                                                                                                                            %          '          V       ^��     �   M   Q   o    �   N   O   o    5�_�                        ����                                                                                                                                                                                                                                                                                                                            4          6          V       ^��     �         r      C   type real_array is array (0 to 15) of integer range -128 to 127;5�_�                        ����                                                                                                                                                                                                                                                                                                                            4          6          V       ^��     �         r      F   type real_Im_array is array (0 to 15) of integer range -128 to 127;5�_�                        ����                                                                                                                                                                                                                                                                                                                            4          6          V       ^��     �                C   type im_array   is array (0 to 15) of integer range -128 to 127;5�_�                        ����                                                                                                                                                                                                                                                                                                                            3          5          V       ^��     �         q      �   constant real_table : real_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);5�_�                        ����                                                                                                                                                                                                                                                                                                                            3          5          V       ^�     �         q      �   constant im_table   : im_array   := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�                    &    ����                                                                                                                                                                                                                                                                                                                            3          5          V       ^�     �         q      �   constant im_table   : real_im_array   := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�                        ����                                                                                                                                                                                                                                                                                                                            3          5          V       ^�     �         q      5   type shiftState is (waitingSvalid, waitingMready);5�_�                        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �         q      8   type axishiftState is (waitingSvalid, waitingMready);5�_�                        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �         q      3   type axiState is (waitingSvalid, waitingMready);5�_�                        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �         q      5   signal state        : shiftState := waitingSvalid;5�_�                         ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ^�$     �                F   type real_im_array is array (0 to 15) of integer range -128 to 127;   �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);   �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�                        ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ^�&     �         n    �         n    5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       ^�-     �                4   type axiStates is (waitingSvalid, waitingMready);5�_�                        ����                                                                                                                                                                                                                                                                                                                                                V       ^�/     �         p    �         p    5�_�                        ����                                                                                                                                                                                                                                                                                                                                                V       ^�0   9 �         q    5�_�                 M        ����                                                                                                                                                                                                                                                                                                                            M           P           V        ^�?     �   o   q   r         end process shift_reg;�   n   p   r            end if;�   m   o   r               end if;�   l   n   r                  end case;�   k   m   r                        end if;�   j   l   r                           end if;�   i   k   r      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   h   j   r      -                        s_axis_tready <= '1';�   g   i   r      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   f   h   r                           else�   e   g   r      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   d   f   r      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   c   e   r      Q                     bitCounter := bitCounter+1;                     --incremento�   b   d   r      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   a   c   r      $               when waitingMready =>�   `   b   r                        end if;�   _   a   r                           state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   ^   `   r      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   ]   _   r      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   \   ^   r      *                     bitCounter      := 0;�   [   ]   r      ,                     s_axis_tready   <= '0';�   Z   \   r      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   Y   [   r      $               when waitingSvalid =>�   X   Z   r                  case state is�   W   Y   r               else�   V   X   r      -            m_axis_tdata  <= (others => '0');�   U   W   r      !            m_axis_tvalid <= '0';�   T   V   r      !            s_axis_tready <= '1';�   S   U   r      +            state         <= waitingSvalid;�   R   T   r               if rst = '0' then�   Q   S   r            if rising_edge(clk) then�   P   R   r         begin�   O   Q   r      <      variable im_part    :std_logic_vector (7    downto 0);�   N   P   r      <      variable real_part  :std_logic_vector (7    downto 0);�   M   O   r      ?      variable index      :integer          range 0      to 15;�   L   N   r      >      variable bitCounter :integer          range 0      to 8;�   K   M   r         mapper_proc:process (clk) is�   I   K   r         end process shift_reg;�   H   J   r            end if;�   G   I   r               end if;�   F   H   r                  end case;�   E   G   r                        end if;�   D   F   r      7                        state         <= waitingSvalid;�   C   E   r      +                        bitCounter    := 0;�   B   D   r      -                        s_axis_tready <= '1';�   A   C   r      -                        m_axis_tvalid <= '0';�   @   B   r      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   r      $               when waitingMready =>�   >   @   r                        end if;�   =   ?   r                           end if;�   <   >   r      7                        state         <= waitingMready;�   ;   =   r      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   r      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   r      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   r      4                     bitCounter   := bitCounter + 1;�   7   9   r                           �   6   8   r      /                     m_axis_tdata <= real_part;�   5   7   r      T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   4   6   r      V                     real_part    := std_logic_vector(to_signed(real_table(index),8));�   3   5   r      T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   r      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   r      $               when waitingSvalid =>�   0   2   r                  case state is�   /   1   r               else�   .   0   r                  bitCounter    := 0;�   -   /   r      -            m_axis_tdata  <= (others => '0');�   ,   .   r      !            m_axis_tvalid <= '0';�   +   -   r      !            s_axis_tready <= '1';�   *   ,   r      +            state         <= waitingSvalid;�   )   +   r               if rst = '0' then�   (   *   r            if rising_edge(clk) then�   '   )   r         begin�   &   (   r      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   r      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   r      ,      variable index :integer range 0 to 15;�   #   %   r      0      variable bitCounter :integer range 0 to 8;�   "   $   r         shift_reg:process (clk) is�          r      4   signal state        : axiStates := waitingSvalid;�         r      4   type axiStates is (waitingSvalid, waitingMready);�         r      �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         r      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         r      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         r      *           rst           : in  STD_LOGIC);�         r      )           clk           : in  STD_LOGIC;�         r      )           s_axis_tready : out STD_LOGIC;�         r      )           s_axis_tlast  : in  STD_LOGIC;�         r      )           s_axis_tvalid : in  STD_LOGIC;�         r      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         r      )           m_axis_tready : in  STD_LOGIC;�   
      r      )           m_axis_tlast  : out STD_LOGIC;�   	      r      )           m_axis_tvalid : out STD_LOGIC;�      
   r      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   r          Port(  �   N   P          8      variable real_part :std_logic_vector (7 downto 0);�   M   O          ,      variable index :integer range 0 to 15;�   L   N          0      variable bitCounter :integer range 0 to 8;�   O   Q          8      variable im_part   :std_logic_vector (7 downto 0);5�_�                 M        ����                                                                                                                                                                                                                                                                                                                            M           P           V        ^�A     �   o   q   r         end process shift_reg;�   n   p   r            end if;�   m   o   r               end if;�   l   n   r                  end case;�   k   m   r                        end if;�   j   l   r                           end if;�   i   k   r      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   h   j   r      -                        s_axis_tready <= '1';�   g   i   r      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   f   h   r                           else�   e   g   r      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   d   f   r      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   c   e   r      Q                     bitCounter := bitCounter+1;                     --incremento�   b   d   r      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   a   c   r      $               when waitingMready =>�   `   b   r                        end if;�   _   a   r                           state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   ^   `   r      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   ]   _   r      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   \   ^   r      *                     bitCounter      := 0;�   [   ]   r      ,                     s_axis_tready   <= '0';�   Z   \   r      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   Y   [   r      $               when waitingSvalid =>�   X   Z   r                  case state is�   W   Y   r               else�   V   X   r      -            m_axis_tdata  <= (others => '0');�   U   W   r      !            m_axis_tvalid <= '0';�   T   V   r      !            s_axis_tready <= '1';�   S   U   r      +            state         <= waitingSvalid;�   R   T   r               if rst = '0' then�   Q   S   r            if rising_edge(clk) then�   P   R   r         begin�   O   Q   r      ?      variable im_part    :std_logic_vector ( 7    downto 0 ) ;�   N   P   r      ?      variable real_part  :std_logic_vector ( 7    downto 0 ) ;�   M   O   r      ?      variable index      :integer          range 0      to 15;�   L   N   r      ?      variable bitCounter :integer          range 0      to 8 ;�   K   M   r         mapper_proc:process (clk) is�   I   K   r         end process shift_reg;�   H   J   r            end if;�   G   I   r               end if;�   F   H   r                  end case;�   E   G   r                        end if;�   D   F   r      7                        state         <= waitingSvalid;�   C   E   r      +                        bitCounter    := 0;�   B   D   r      -                        s_axis_tready <= '1';�   A   C   r      -                        m_axis_tvalid <= '0';�   @   B   r      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   r      $               when waitingMready =>�   >   @   r                        end if;�   =   ?   r                           end if;�   <   >   r      7                        state         <= waitingMready;�   ;   =   r      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   r      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   r      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   r      4                     bitCounter   := bitCounter + 1;�   7   9   r                           �   6   8   r      /                     m_axis_tdata <= real_part;�   5   7   r      T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   4   6   r      V                     real_part    := std_logic_vector(to_signed(real_table(index),8));�   3   5   r      T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   r      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   r      $               when waitingSvalid =>�   0   2   r                  case state is�   /   1   r               else�   .   0   r                  bitCounter    := 0;�   -   /   r      -            m_axis_tdata  <= (others => '0');�   ,   .   r      !            m_axis_tvalid <= '0';�   +   -   r      !            s_axis_tready <= '1';�   *   ,   r      +            state         <= waitingSvalid;�   )   +   r               if rst = '0' then�   (   *   r            if rising_edge(clk) then�   '   )   r         begin�   &   (   r      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   r      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   r      ,      variable index :integer range 0 to 15;�   #   %   r      0      variable bitCounter :integer range 0 to 8;�   "   $   r         shift_reg:process (clk) is�          r      4   signal state        : axiStates := waitingSvalid;�         r      4   type axiStates is (waitingSvalid, waitingMready);�         r      �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         r      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         r      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         r      *           rst           : in  STD_LOGIC);�         r      )           clk           : in  STD_LOGIC;�         r      )           s_axis_tready : out STD_LOGIC;�         r      )           s_axis_tlast  : in  STD_LOGIC;�         r      )           s_axis_tvalid : in  STD_LOGIC;�         r      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         r      )           m_axis_tready : in  STD_LOGIC;�   
      r      )           m_axis_tlast  : out STD_LOGIC;�   	      r      )           m_axis_tvalid : out STD_LOGIC;�      
   r      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   r          Port(  �   N   P          <      variable real_part  :std_logic_vector (7    downto 0);�   M   O          ?      variable index      :integer          range 0      to 15;�   L   N          >      variable bitCounter :integer          range 0      to 8;�   O   Q          <      variable im_part    :std_logic_vector (7    downto 0);5�_�                 M   #    ����                                                                                                                                                                                                                                                                                                                            M   #       N   +          +    ^�F     �   L   O   r      ?      variable bitCounter :integer          range 0      to 8 ;   ?      variable index      :integer          range 0      to 15;5�_�                 M   +    ����                                                                                                                                                                                                                                                                                                                            M   +       N   /          /    ^�I     �   L   O   r      6      variable bitCounter :integer range 0      to 8 ;   6      variable index      :integer range 0      to 15;5�_�                  O   0    ����                                                                                                                                                                                                                                                                                                                            O   0       P   2          2    ^�K     �   N   Q   r      ?      variable real_part  :std_logic_vector ( 7    downto 0 ) ;   ?      variable im_part    :std_logic_vector ( 7    downto 0 ) ;5�_�    !              ^        ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�n     �   ]   b   r    �   ^   _   r    5�_�     "          !   a       ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�r     �   a   c   v    5�_�  !  #          "   c       ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�v     �   b   c          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�  "  %          #   b        ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�w     �   a   b           5�_�  #  &  $      %   ^        ����                                                                                                                                                                                                                                                                                                                            ^          c          V       ^�}     �   r   t   u         end process shift_reg;�   q   s   u            end if;�   p   r   u               end if;�   o   q   u                  end case;�   n   p   u                        end if;�   m   o   u                           end if;�   l   n   u      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   k   m   u      -                        s_axis_tready <= '1';�   j   l   u      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   i   k   u                           else�   h   j   u      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   g   i   u      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   f   h   u      Q                     bitCounter := bitCounter+1;                     --incremento�   e   g   u      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   d   f   u      $               when waitingMready =>�   c   e   u                        end if;�   b   d   u      }                     state         <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   a   c   u      o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   `   b   u      0                     m_axis_tdata  <= real_part;�   _   a   u      U                     im_part       := std_logic_vector(to_signed(im_table(index),8));�   ^   `   u      W                     real_part     := std_logic_vector(to_signed(real_table(index),8));�   ]   _   u      U                     index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   \   ^   u      *                     bitCounter      := 0;�   [   ]   u      ,                     s_axis_tready   <= '0';�   Z   \   u      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   Y   [   u      $               when waitingSvalid =>�   X   Z   u                  case state is�   W   Y   u               else�   V   X   u      -            m_axis_tdata  <= (others => '0');�   U   W   u      !            m_axis_tvalid <= '0';�   T   V   u      !            s_axis_tready <= '1';�   S   U   u      +            state         <= waitingSvalid;�   R   T   u               if rst = '0' then�   Q   S   u            if rising_edge(clk) then�   P   R   u         begin�   O   Q   u      <      variable im_part    :std_logic_vector ( 7 downto 0 ) ;�   N   P   u      <      variable real_part  :std_logic_vector ( 7 downto 0 ) ;�   M   O   u      1      variable index      :integer range 0 to 15;�   L   N   u      1      variable bitCounter :integer range 0 to 8 ;�   K   M   u         mapper_proc:process (clk) is�   I   K   u         end process shift_reg;�   H   J   u            end if;�   G   I   u               end if;�   F   H   u                  end case;�   E   G   u                        end if;�   D   F   u      7                        state         <= waitingSvalid;�   C   E   u      +                        bitCounter    := 0;�   B   D   u      -                        s_axis_tready <= '1';�   A   C   u      -                        m_axis_tvalid <= '0';�   @   B   u      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   u      $               when waitingMready =>�   >   @   u                        end if;�   =   ?   u                           end if;�   <   >   u      7                        state         <= waitingMready;�   ;   =   u      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   u      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   u      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   u      4                     bitCounter   := bitCounter + 1;�   7   9   u                           �   6   8   u      /                     m_axis_tdata <= real_part;�   5   7   u      T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   4   6   u      V                     real_part    := std_logic_vector(to_signed(real_table(index),8));�   3   5   u      T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   u      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   u      $               when waitingSvalid =>�   0   2   u                  case state is�   /   1   u               else�   .   0   u                  bitCounter    := 0;�   -   /   u      -            m_axis_tdata  <= (others => '0');�   ,   .   u      !            m_axis_tvalid <= '0';�   +   -   u      !            s_axis_tready <= '1';�   *   ,   u      +            state         <= waitingSvalid;�   )   +   u               if rst = '0' then�   (   *   u            if rising_edge(clk) then�   '   )   u         begin�   &   (   u      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   u      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   u      ,      variable index :integer range 0 to 15;�   #   %   u      0      variable bitCounter :integer range 0 to 8;�   "   $   u         shift_reg:process (clk) is�          u      4   signal state        : axiStates := waitingSvalid;�         u      4   type axiStates is (waitingSvalid, waitingMready);�         u      �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         u      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         u      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         u      *           rst           : in  STD_LOGIC);�         u      )           clk           : in  STD_LOGIC;�         u      )           s_axis_tready : out STD_LOGIC;�         u      )           s_axis_tlast  : in  STD_LOGIC;�         u      )           s_axis_tvalid : in  STD_LOGIC;�         u      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         u      )           m_axis_tready : in  STD_LOGIC;�   
      u      )           m_axis_tlast  : out STD_LOGIC;�   	      u      )           m_axis_tvalid : out STD_LOGIC;�      
   u      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   u          Port(  �   ]   _          T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   b   d                               state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   a   c          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   `   b          /                     m_axis_tdata <= real_part;�   _   a          T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   ^   `          V                     real_part    := std_logic_vector(to_signed(real_table(index),8));5�_�  %  '          &   \        ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   r   t   u         end process shift_reg;�   q   s   u            end if;�   p   r   u               end if;�   o   q   u                  end case;�   n   p   u                        end if;�   m   o   u                           end if;�   l   n   u      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   k   m   u      -                        s_axis_tready <= '1';�   j   l   u      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   i   k   u                           else�   h   j   u      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   g   i   u      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   f   h   u      Q                     bitCounter := bitCounter+1;                     --incremento�   e   g   u      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   d   f   u      $               when waitingMready =>�   c   e   u                        end if;�   b   d   u      }                     state         <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   a   c   u      o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   `   b   u      0                     m_axis_tdata  <= real_part;�   _   a   u      U                     im_part       := std_logic_vector(to_signed(im_table(index),8));�   ^   `   u      W                     real_part     := std_logic_vector(to_signed(real_table(index),8));�   ]   _   u      U                     index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   \   ^   u      (                     bitCounter    := 0;�   [   ]   u      *                     s_axis_tready <= '0';�   Z   \   u      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   Y   [   u      $               when waitingSvalid =>�   X   Z   u                  case state is�   W   Y   u               else�   V   X   u      -            m_axis_tdata  <= (others => '0');�   U   W   u      !            m_axis_tvalid <= '0';�   T   V   u      !            s_axis_tready <= '1';�   S   U   u      +            state         <= waitingSvalid;�   R   T   u               if rst = '0' then�   Q   S   u            if rising_edge(clk) then�   P   R   u         begin�   O   Q   u      <      variable im_part    :std_logic_vector ( 7 downto 0 ) ;�   N   P   u      <      variable real_part  :std_logic_vector ( 7 downto 0 ) ;�   M   O   u      1      variable index      :integer range 0 to 15;�   L   N   u      1      variable bitCounter :integer range 0 to 8 ;�   K   M   u         mapper_proc:process (clk) is�   I   K   u         end process shift_reg;�   H   J   u            end if;�   G   I   u               end if;�   F   H   u                  end case;�   E   G   u                        end if;�   D   F   u      7                        state         <= waitingSvalid;�   C   E   u      +                        bitCounter    := 0;�   B   D   u      -                        s_axis_tready <= '1';�   A   C   u      -                        m_axis_tvalid <= '0';�   @   B   u      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   ?   A   u      $               when waitingMready =>�   >   @   u                        end if;�   =   ?   u                           end if;�   <   >   u      7                        state         <= waitingMready;�   ;   =   u      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   :   <   u      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   9   ;   u      \                     if bitCounter = 1 then                             --porque bit voy?   �   8   :   u      4                     bitCounter   := bitCounter + 1;�   7   9   u                           �   6   8   u      /                     m_axis_tdata <= real_part;�   5   7   u      T                     im_part      := std_logic_vector(to_signed(im_table(index),8));�   4   6   u      V                     real_part    := std_logic_vector(to_signed(real_table(index),8));�   3   5   u      T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   2   4   u      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   1   3   u      $               when waitingSvalid =>�   0   2   u                  case state is�   /   1   u               else�   .   0   u                  bitCounter    := 0;�   -   /   u      -            m_axis_tdata  <= (others => '0');�   ,   .   u      !            m_axis_tvalid <= '0';�   +   -   u      !            s_axis_tready <= '1';�   *   ,   u      +            state         <= waitingSvalid;�   )   +   u               if rst = '0' then�   (   *   u            if rising_edge(clk) then�   '   )   u         begin�   &   (   u      8      variable im_part   :std_logic_vector (7 downto 0);�   %   '   u      8      variable real_part :std_logic_vector (7 downto 0);�   $   &   u      ,      variable index :integer range 0 to 15;�   #   %   u      0      variable bitCounter :integer range 0 to 8;�   "   $   u         shift_reg:process (clk) is�          u      4   signal state        : axiStates := waitingSvalid;�         u      4   type axiStates is (waitingSvalid, waitingMready);�         u      �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         u      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         u      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         u      *           rst           : in  STD_LOGIC);�         u      )           clk           : in  STD_LOGIC;�         u      )           s_axis_tready : out STD_LOGIC;�         u      )           s_axis_tlast  : in  STD_LOGIC;�         u      )           s_axis_tvalid : in  STD_LOGIC;�         u      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         u      )           m_axis_tready : in  STD_LOGIC;�   
      u      )           m_axis_tlast  : out STD_LOGIC;�   	      u      )           m_axis_tvalid : out STD_LOGIC;�      
   u      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   u          Port(  �   [   ]          ,                     s_axis_tready   <= '0';�   b   d          }                     state         <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   a   c          o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   `   b          0                     m_axis_tdata  <= real_part;�   _   a          U                     im_part       := std_logic_vector(to_signed(im_table(index),8));�   ^   `          W                     real_part     := std_logic_vector(to_signed(real_table(index),8));�   ]   _          U                     index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));�   \   ^          *                     bitCounter      := 0;5�_�  &  (          '   h   #    ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   g   i   u      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�  '  )          (   h   %    ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   g   i   u      f                     if bitCounter = 8 then                             --perfecto, porque bit voy?   5�_�  (  *          )   h   #    ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   g   i   u      f                     if bitCounter = 1 then                             --perfecto, porque bit voy?   5�_�  )  +          *   h   %    ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   g   i   u      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   5�_�  *  ,          +   i   %    ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   h   j   u    �   i   j   u    5�_�  +  .          ,   i       ����                                                                                                                                                                                                                                                                                                                            \           c           V        ^��     �   h   j          0                     m_axis_tdata  <= real_part;5�_�  ,  /  -      .   i   )    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^��     �   h   j   v      3                        m_axis_tdata  <= real_part;5�_�  .  0          /   j       ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^��     �   i   j          W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�  /  1          0   s       ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^��     �   r   t   u         end process shift_reg;5�_�  0  2          1   f   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   e   g   u      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�  1  3          2   f   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   e   g   u      p                  if m_axis_tready = '1' then                          --lo puedo empezar a mandar al otro lado?5�_�  2  4          3   f   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   e   g   u      o                  if m_axis_tready = '1' then                         --lo puedo empezar a mandar al otro lado?5�_�  3  5          4   f   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   e   g   u      n                  if m_axis_tready = '1' then                        --lo puedo empezar a mandar al otro lado?5�_�  4  6          5   f   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   e   g   u      m                  if m_axis_tready = '1' then                       --lo puedo empezar a mandar al otro lado?5�_�  5  7          6   g   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   f   h   u      Q                     bitCounter := bitCounter+1;                     --incremento5�_�  6  8          7   g   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   f   h   u      P                     bitCounter := bitCounter+1;                    --incremento5�_�  7  9          8   h   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   g   i   u      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   5�_�  8  :          9   h   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   g   i   u      e                     if bitCounter < 2 then                            --perfecto, porque bit voy?   5�_�  9  ;          :   h   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   g   i   u      d                     if bitCounter < 2 then                           --perfecto, porque bit voy?   5�_�  :  <          ;   h   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   g   i   u      c                     if bitCounter < 2 then                          --perfecto, porque bit voy?   5�_�  ;  =          <   h   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   g   i   u      b                     if bitCounter < 2 then                         --perfecto, porque bit voy?   5�_�  <  >          =   k   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   j   l   u      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  =  ?          >   k   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   j   l   u      �                        m_axis_tvalid <= '0' ;                         --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  >  @          ?   k   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   j   l   u      �                        m_axis_tvalid <= '0' ;                        --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  ?  A          @   k   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   j   l   u      �                        m_axis_tvalid <= '0' ;                       --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  @  B          A   k   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   j   l   u      �                        m_axis_tvalid <= '0' ;                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  A  C          B   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�  B  D          C   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;                   --cambio de estado, y le doy un clk para que ponga el dato5�_�  C  E          D   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;                  --cambio de estado, y le doy un clk para que ponga el dato5�_�  D  F          E   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;                 --cambio de estado, y le doy un clk para que ponga el dato5�_�  E  G          F   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;                --cambio de estado, y le doy un clk para que ponga el dato5�_�  F  H          G   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      �                        state         <= waitingSvalid;               --cambio de estado, y le doy un clk para que ponga el dato5�_�  G  I          H   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u                              state         <= waitingSvalid;              --cambio de estado, y le doy un clk para que ponga el dato5�_�  H  J          I   m   C    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^�     �   l   n   u      ~                        state         <= waitingSvalid;             --cambio de estado, y le doy un clk para que ponga el dato5�_�  I  K          J   #       ����                                                                                                                                                                                                                                                                                                                            J          #          V   C    ^�     �   "   #       (      shift_reg:process (clk) is   0      variable bitCounter :integer range 0 to 8;   ,      variable index :integer range 0 to 15;   8      variable real_part :std_logic_vector (7 downto 0);   8      variable im_part   :std_logic_vector (7 downto 0);      begin         if rising_edge(clk) then            if rst = '0' then   +            state         <= waitingSvalid;   !            s_axis_tready <= '1';   !            m_axis_tvalid <= '0';   -            m_axis_tdata  <= (others => '0');               bitCounter    := 0;            else               case state is   $               when waitingSvalid =>   r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   T                     index        := to_integer(unsigned(s_axis_tdata(3 downto 0)));   V                     real_part    := std_logic_vector(to_signed(real_table(index),8));   T                     im_part      := std_logic_vector(to_signed(im_table(index),8));   /                     m_axis_tdata <= real_part;                           4                     bitCounter   := bitCounter + 1;   \                     if bitCounter = 1 then                             --porque bit voy?      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo   `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada   7                        state         <= waitingMready;                        end if;                     end if;   $               when waitingMready =>   �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..   -                        m_axis_tvalid <= '0';   -                        s_axis_tready <= '1';   +                        bitCounter    := 0;   7                        state         <= waitingSvalid;                     end if;               end case;            end if;         end if;      end process shift_reg;5�_�  J  L          K   #        ����                                                                                                                                                                                                                                                                                                                            #          #          V   C    ^�     �   "   #           5�_�  K  M          L   "        ����                                                                                                                                                                                                                                                                                                                            #          #          V   C    ^�     �   !   "           5�_�  L  N          M           ����                                                                                                                                                                                                                                                                                                                                                  V       ^�     �                     5�_�  M  O          N           ����                                                                                                                                                                                                                                                                                                                                                  V       ^�     �                W--junto 8 bytes en uno, tomando solo el bit 0 de cada byte y lo mando por el axi master5�_�  N  P          O           ����                                                                                                                                                                                                                                                                                                                                                  V       ^�   : �                 5�_�  O  Q          P   ,        ����                                                                                                                                                                                                                                                                                                                                                             ^/J     �   +   6   G    �   ,   -   G    5�_�  P  S          Q   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^/O     �   +   -   Q    �   ,   -   Q    5�_�  Q  T  R      S   0   @    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   /   1   R      B                     bitCounter                 := bitCounter + 2;5�_�  S  U          T   .   3    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   -   /   R      C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);5�_�  T  V          U   1   %    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   0   2   R      \                     if bitCounter = 8 then                             --porque bit voy?   5�_�  U  W          V   1   #    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   0   2   R      \                     if bitCounter = 1 then                             --porque bit voy?   5�_�  V  X          W   1   %    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   0   2   R      \                     if bitCounter < 1 then                             --porque bit voy?   5�_�  W  Y          X   1   #    ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   0   2   R      \                     if bitCounter < 2 then                             --porque bit voy?   5�_�  X  Z          Y   .   "    ����                                                                                                                                                                                                                                                                                                                            .   "       /   "          "    ^/�     �   .   0   R      C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);�   -   /   R      C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);5�_�  Y  [          Z   .   "    ����                                                                                                                                                                                                                                                                                                                            .   "       /   #          #    ^0�     �   -   0   R      E                     m_axis_tdata(4-bitCounter)   <= s_axis_tdata(0);   E                     m_axis_tdata(4-bitCounter+1) <= s_axis_tdata(1);5�_�  Z  \          [   0   @    ����                                                                                                                                                                                                                                                                                                                            .   "       /   #          #    ^0�     �   /   1   R      B                     bitCounter                 := bitCounter + 1;5�_�  [  ]          \   1   %    ����                                                                                                                                                                                                                                                                                                                            .   "       /   #          #    ^0�     �   0   2   R      \                     if bitCounter = 2 then                             --porque bit voy?   5�_�  \  ^          ]   "   %    ����                                                                                                                                                                                                                                                                                                                            .   "       /   #          #    ^1D     �   !   #   R    �   "   #   R    5�_�  ]  _          ^   #       ����                                                                                                                                                                                                                                                                                                                            /   "       0   #          #    ^1G     �   "   $   S      <      variable im_part    :std_logic_vector ( 7 downto 0 ) ;5�_�  ^  `          _   #       ����                                                                                                                                                                                                                                                                                                                            /   "       0   #          #    ^1K     �   "   $   S      =      variable data2Map    :std_logic_vector ( 7 downto 0 ) ;5�_�  _  a          `   #   .    ����                                                                                                                                                                                                                                                                                                                            /   "       0   #          #    ^1P     �   "   $   S      <      variable data2Map   :std_logic_vector ( 7 downto 0 ) ;5�_�  `  b          a   #   .    ����                                                                                                                                                                                                                                                                                                                            /   "       0   #          #    ^1R     �   "   $   S      <      variable data2Map   :std_logic_vector ( 4 downto 0 ) ;5�_�  a  c          b   /       ����                                                                                                                                                                                                                                                                                                                            /          0                 ^1Y     �   .   1   S      C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);   C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);5�_�  b  d          c   /       ����                                                                                                                                                                                                                                                                                                                            /          0                   ^1`     �   .   0   S      7                     (bitCounter)   <= s_axis_tdata(0);�   .   1   S      C                     e_axis_tdata(bitCounter)   <= s_axis_tdata(0);   C                     e_axis_tdata(bitCounter+1) <= s_axis_tdata(1);5�_�  c  e          d   3        ����                                                                                                                                                                                                                                                                                                                            <          =          V       ^1z     �   2   5   S    �   3   4   S    5�_�  d  f          e   3        ����                                                                                                                                                                                                                                                                                                                            3          4          V       ^1|     �   3   5          W                     real_part     := std_logic_vector(to_signed(real_table(index),8));�   2   4          U                     index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));5�_�  e  g          f   3   =    ����                                                                                                                                                                                                                                                                                                                            3          4          V       ^1�     �   2   4   U      X                        index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));5�_�  f  h          g   3   E    ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   2   4   U      T                        index         := to_integer(unsigned(data2Map(3 downto 0)));5�_�  g  i          h   4       ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   3   5   U      Z                        real_part     := std_logic_vector(to_signed(real_table(index),8));5�_�  h  j          i   4   %    ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   3   5   U      ]                        m_axis_tdata     := std_logic_vector(to_signed(real_table(index),8));5�_�  i  k          j   4   %    ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   3   5   U      \                        m_axis_tdata    := std_logic_vector(to_signed(real_table(index),8));5�_�  j  l          k   4   %    ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   3   5   U      [                        m_axis_tdata   := std_logic_vector(to_signed(real_table(index),8));5�_�  k  m          l   4   &    ����                                                                                                                                                                                                                                                                                                                            3   E       3   P       v   P    ^1�     �   3   5   U      Z                        m_axis_tdata  := std_logic_vector(to_signed(real_table(index),8));5�_�  l  n          m   1   ,    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   0   2   U      B                     bitCounter                 := bitCounter + 2;5�_�  m  o          n   7   ,    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   6   8   U    �   7   8   U    5�_�  n  p          o   7       ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   6   8   V      >                     bitCounter             := bitCounter + 2;5�_�  o  q          p   7   &    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   6   8   V      A                        bitCounter             := bitCounter + 2;5�_�  p  r          q   7   )    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   6   8   V      8                        bitCounter    := bitCounter + 2;5�_�  q  s          r   7   )    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^1�     �   6   8   V      *                        bitCounter    := ;5�_�  r  t          s   J   $    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^2     �   I   K   V    �   J   K   V    5�_�  s  u          t   J   D    ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^2     �   I   K   W      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));5�_�  t  v          u   K       ����                                                                                                                                                                                                                                                                                                                            1   &       /   &       V   &    ^2     �   J   K          1                        m_axis_tdata  <= im_part;5�_�  u  w          v   ;       ����                                                                                                                                                                                                                                                                                                                            E          ;          V       ^2#     �   :   ;          $               when waitingSvalid =>   r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   *                     s_axis_tready <= '0';   (                     bitCounter    := 0;   U                     index         := to_integer(unsigned(s_axis_tdata(3 downto 0)));   W                     real_part     := std_logic_vector(to_signed(real_table(index),8));   U                     im_part       := std_logic_vector(to_signed(im_table(index),8));   0                     m_axis_tdata  <= real_part;   o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato   }                     state         <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato                     end if;5�_�  v  x          w   !        ����                                                                                                                                                                                                                                                                                                                            !          "          V       ^2:     �       !          <      variable real_part  :std_logic_vector ( 7 downto 0 ) ;   <      variable im_part    :std_logic_vector ( 7 downto 0 ) ;5�_�  w  y          x   A       ����                                                                                                                                                                                                                                                                                                                            !          !          V       ^2]   = �   @   B   I    �   A   B   I    5�_�  x  z          y   !       ����                                                                                                                                                                                                                                                                                                                                                             ^6     �       "   J      <      variable data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  y  {          z   !       ����                                                                                                                                                                                                                                                                                                                                                             ^6   > �       "   J      :      signal data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  z  |          {   !        ����                                                                                                                                                                                                                                                                                                                            !          !          V       ^6     �       !          <      signal   data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  {  }          |           ����                                                                                                                                                                                                                                                                                                                            !          !          V       ^6     �         I    �         I    5�_�  |  ~          }          ����                                                                                                                                                                                                                                                                                                                            "          "          V       ^6     �                <      signal   data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  }            ~      
    ����                                                                                                                                                                                                                                                                                                                            "          "          V       ^6      �         J      9   signal   data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  ~  �                
    ����                                                                                                                                                                                                                                                                                                                            "          "          V       ^6"     �         J      8   signal  data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�    �          �          ����                                                                                                                                                                                                                                                                                                                            "          "          V       ^6$   @ �         J      4   signal state        : axiStates := waitingSvalid;5�_�  �  �  �      �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^9M   A �         J      end mapper;�         J      entity mapper is5�_�  �  �  �      �   #       ����                                                                                                                                                                                                                                                                                                                            #          G                 ^�7   B �   #   H   J   $            if rst = '0' then   +            state         <= waitingSvalid;   !            s_axis_tready <= '1';   !            m_axis_tvalid <= '0';   -            m_axis_tdata  <= (others => '0');            else               case state is   $               when waitingSvalid =>   r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   ?                     data2Map(bitCounter)   <= s_axis_tdata(0);   ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);   >                     bitCounter             := bitCounter + 2;   \                     if bitCounter = 4 then                             --porque bit voy?      H                        index         := to_integer(unsigned(data2Map));   Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo   `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada   +                        bitCounter    := 0;   7                        state         <= waitingMready;                        end if;                     end if;   $               when waitingMready =>   l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   O                     bitCounter := bitCounter+1;                   --incremento   a                     if bitCounter < 2 then                        --perfecto, porque bit voy?      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));                        else   �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   -                        s_axis_tready <= '1';   +                        bitCounter    := 0;   }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato                        end if;                     end if;               end case;            end if;         end if;�   "   $   J            if rising_edge(clk) then5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�E     �   "   9   J             --if rising_edge(clk) then         --   if rst = '0' then   -      --      state         <= waitingSvalid;   #      --      s_axis_tready <= '1';   #      --      m_axis_tvalid <= '0';   /      --      m_axis_tdata  <= (others => '0');         --   else         --      case state is   &      --         when waitingSvalid =>   t      --            if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   A      --               data2Map(bitCounter)   <= s_axis_tdata(0);   A      --               data2Map(bitCounter+1) <= s_axis_tdata(1);   @      --               bitCounter             := bitCounter + 2;   ^      --               if bitCounter = 4 then                             --porque bit voy?      J      --                  index         := to_integer(unsigned(data2Map));   \      --                  m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   n      --                  s_axis_tready <= '0';                              --entonces yo tambien estoy listo   b      --                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada   -      --                  bitCounter    := 0;   9      --                  state         <= waitingMready;         --               end if;         --            end if;5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�J     �   F   H   J            --end if;5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�J     �   F   H   J            -end if;5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�P     �   D   F   J            --      end case;5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�P     �   D   F   J            -      end case;5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�Q     �   E   G   J            --   end if;5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�Q   D �   E   G   J            -   end if;5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�h     �   8   :   J      &      --         when waitingMready =>5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�h     �   8   :   J      %      -         when waitingMready =>5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�n     �   D   F   J    �   E   F   J    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            #          8                 ^�o   E �   D   F   K      $               when waitingMready =>5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                            0          7                 ^��   F �   0   8   K      H                        index         := to_integer(unsigned(data2Map));   Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo   `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada   +                        bitCounter    := 0;   7                        state         <= waitingMready;                        end if;�   /   1   K      \                     if bitCounter = 4 then                             --porque bit voy?   5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                            0          7                 ^��     �   /   1   K      ^                     --if bitCounter = 4 then                             --porque bit voy?   5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                            0          7                 ^��     �   /   1   K      ]                     -if bitCounter = 4 then                             --porque bit voy?   5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                            0          7                 ^��     �   6   8   K                           --end if;5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                            0          7                 ^��   G �   6   8   K                           -end if;5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          6                 ^��     �   0   7   K      J                     --   index         := to_integer(unsigned(data2Map));   \                     --   m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   n                     --   s_axis_tready <= '0';                              --entonces yo tambien estoy listo   b                     --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada   -                     --   bitCounter    := 0;   9                     --   state         <= waitingMready;5�_�  �  �          �   1        ����                                                                                                                                                                                                                                                                                                                            1          6          V       ^��   K �   5   7          6                       state         <= waitingMready;�   4   6          *                       bitCounter    := 0;�   3   5          _                       m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   2   4          k                       s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   1   3          Y                       m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   0   2          G                       index         := to_integer(unsigned(data2Map));5�_�  �  �  �      �   :       ����                                                                                                                                                                                                                                                                                                                            :          D                 ^��   L �   9   E   K      n      --            if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   Q      --               bitCounter := bitCounter+1;                   --incremento   c      --               if bitCounter < 2 then                        --perfecto, porque bit voy?      Z      --                  m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));         --               else   �      --                  m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   /      --                  s_axis_tready <= '1';   -      --                  bitCounter    := 0;         --                  state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato         --               end if;         --            end if;5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            :          D                 ^�     �   0   2   K      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            :          D                 ^�     �   1   3   K    �   2   3   K    5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�     �   1   3   L      J                        --index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�     �   1   3   L      I                        -index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2   )    ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�     �   1   3   L      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2   )    ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�   N �   1   3   L      )                        index         := 5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�     �   0   2   L      J                        --index         := to_integer(unsigned(data2Map));5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�     �   0   2   L      I                        -index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            ;          E                 ^�    Q �   1   2          +                        index         := 0;5�_�  �  �  �      �      )    ����                                                                                                                                                                                                                                                                                                                            :          D                 ^��   R �         K      7   signal data2Map   :std_logic_vector ( 3 downto 0 ) ;5�_�  �  �          �   !   )    ����                                                                                                                                                                                                                                                                                                                            :          D                 ^��   S �       "   K      1      variable index      :integer range 0 to 15;5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            :          D                 ^��     �       "   K      3      variable index      :integer range -16 to 15;5�_�  �  �          �   !   )    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��   T �       "   K      3      variable index      :natural range -16 to 15;5�_�  �  �  �      �           ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�g   V �      !   K      1      variable bitCounter :integer range 0 to 8 ;5�_�  �  �  �      �   1       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   0   2   K      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   1   3   K    �   2   3   K    5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   1   3   L      J                        --index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   1   3   L      I                        -index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2   )    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   1   3   L      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2   )    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��   X �   1   3   L      )                        index         := 5�_�  �  �  �      �   (       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�*     �   '   )   L    �   (   )   L    5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�+     �   (   *   M      -            m_axis_tdata  <= (others => '0');5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�1     �   (   *   M      )            data2Map  <= (others => '0');5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�2   Y �   (   *   M      )            data2Map  "= (others => '0');5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�C     �   (   *   M      )            data2Map  := (others => '0');5�_�  �  �          �   %        ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�F   Z �   J   L   M         end process mapper_proc;�   I   K   M            end if;�   H   J   M               end if;�   G   I   M                  end case;�   F   H   M                     when others =>�   E   G   M                        end if;�   D   F   M                           end if;�   C   E   M      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   B   D   M      +                        bitCounter    := 0;�   A   C   M      -                        s_axis_tready <= '1';�   @   B   M      �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   ?   A   M                           else�   >   @   M      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));�   =   ?   M      a                     if bitCounter < 2 then                        --perfecto, porque bit voy?   �   <   >   M      O                     bitCounter := bitCounter+1;                   --incremento�   ;   =   M      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   :   <   M      $               when waitingMready =>�   9   ;   M                        end if;�   8   :   M                           end if;�   7   9   M      7                        state         <= waitingMready;�   6   8   M      +                        bitCounter    := 0;�   5   7   M      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   4   6   M      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   3   5   M      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   2   4   M      +                        index         := 0;�   1   3   M      J                        --index         := to_integer(unsigned(data2Map));�   0   2   M      \                     if bitCounter = 4 then                             --porque bit voy?   �   /   1   M      >                     bitCounter             := bitCounter + 2;�   .   0   M      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   -   /   M      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   ,   .   M      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   +   -   M      $               when waitingSvalid =>�   *   ,   M                  case state is�   )   +   M               else�   (   *   M      -            data2Map      <= (others => '0');�   '   )   M      -            m_axis_tdata  <= (others => '0');�   &   (   M      !            m_axis_tvalid <= '0';�   %   '   M      !            s_axis_tready <= '1';�   $   &   M      +            state         <= waitingSvalid;�   #   %   M               if rst = '0' then�   "   $   M            if rising_edge(clk) then�   !   #   M         begin�       "   M      1      variable index      :natural range 0 to 15;�      !   M      1      variable bitCounter :natural range 0 to 8 ;�          M         mapper_proc:process (clk) is�         M      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;�         M      2   signal state      : axiStates := waitingSvalid;�         M      4   type axiStates is (waitingSvalid, waitingMready);�         M      �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         M      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         M      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         M      *           rst           : in  STD_LOGIC);�         M      )           clk           : in  STD_LOGIC;�         M      )           s_axis_tready : out STD_LOGIC;�         M      )           s_axis_tlast  : in  STD_LOGIC;�         M      )           s_axis_tvalid : in  STD_LOGIC;�         M      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   	      M      )           m_axis_tready : in  STD_LOGIC;�      
   M      )           m_axis_tlast  : out STD_LOGIC;�      	   M      )           m_axis_tvalid : out STD_LOGIC;�         M      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         M          Port(  �   $   &          +            state         <= waitingSvalid;�   &   (          !            m_axis_tvalid <= '0';�   %   '          !            s_axis_tready <= '1';�   (   *          )            data2Map  <= (others => '0');�   '   )          -            m_axis_tdata  <= (others => '0');5�_�  �  �  �      �   2       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�P     �   1   3   M      J                        --index         := to_integer(unsigned(data2Map));5�_�  �  �  �      �   2       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^��   ` �   1   3   M      I                        -index         := to_integer(unsigned(data2Map));5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^��   a �   2   4   M      +                        index         := 0;5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^��   b �   2   3          -                        --index         := 0;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                       J           V        ^��   c �   I   K   L         end process mapper_proc;�          L         mapper_proc:process (clk) is5�_�  �  �  �      �           ����                                                                                                                                                                                                                                                                                                                               �          �       V   �    ^L�     �   I   K   L      !   end process mapper_proc; --}}}�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L                     when others =>�   D   F   L                        end if;�   C   E   L                           end if;�   B   D   L      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   A   C   L      +                        bitCounter    := 0;�   @   B   L      -                        s_axis_tready <= '1';�   ?   A   L      �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   >   @   L                           else�   =   ?   L      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));�   <   >   L      a                     if bitCounter < 2 then                        --perfecto, porque bit voy?   �   ;   =   L      O                     bitCounter := bitCounter+1;                   --incremento�   :   <   L      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   9   ;   L      $               when waitingMready =>�   8   :   L                        end if;�   7   9   L                           end if;�   6   8   L      7                        state         <= waitingMready;�   5   7   L      +                        bitCounter    := 0;�   4   6   L      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   3   5   L      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   2   4   L      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   1   3   L      H                        index         := to_integer(unsigned(data2Map));�   0   2   L      \                     if bitCounter = 4 then                             --porque bit voy?   �   /   1   L      >                     bitCounter             := bitCounter + 2;�   .   0   L      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   -   /   L      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   ,   .   L      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   +   -   L      $               when waitingSvalid =>�   *   ,   L                  case state is�   )   +   L               else�   (   *   L      -            data2Map      <= (others => '0');�   '   )   L      -            m_axis_tdata  <= (others => '0');�   &   (   L      !            m_axis_tvalid <= '0';�   %   '   L      !            s_axis_tready <= '1';�   $   &   L      +            state         <= waitingSvalid;�   #   %   L               if rst = '0' then�   "   $   L            if rising_edge(clk) then�   !   #   L         begin�       "   L      1      variable index      :natural range 0 to 15;�      !   L      1      variable bitCounter :natural range 0 to 8 ;�          L      %   mapper_proc:process (clk) is --{{{�         L      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;�         L      2   signal state      : axiStates := waitingSvalid;�         L      4   type axiStates is (waitingSvalid, waitingMready);�         L      �   constant im_table   : real_im_array  := (25 ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         L      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         L      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         L      *           rst           : in  STD_LOGIC);�         L      )           clk           : in  STD_LOGIC;�         L      )           s_axis_tready : out STD_LOGIC;�         L      )           s_axis_tlast  : in  STD_LOGIC;�         L      )           s_axis_tvalid : in  STD_LOGIC;�         L      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   	      L      )           m_axis_tready : in  STD_LOGIC;�      
   L      )           m_axis_tlast  : out STD_LOGIC;�      	   L      )           m_axis_tvalid : out STD_LOGIC;�         L      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         L          Port(  �                �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�                �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^L�     �   I   K   L      !   end process mapper_proc; --}}}�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L                     when others =>�   D   F   L                        end if;�   C   E   L                           end if;�   B   D   L      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   A   C   L      +                        bitCounter    := 0;�   @   B   L      -                        s_axis_tready <= '1';�   ?   A   L      �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   >   @   L                           else�   =   ?   L      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));�   <   >   L      a                     if bitCounter < 2 then                        --perfecto, porque bit voy?   �   ;   =   L      O                     bitCounter := bitCounter+1;                   --incremento�   :   <   L      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   9   ;   L      $               when waitingMready =>�   8   :   L                        end if;�   7   9   L                           end if;�   6   8   L      7                        state         <= waitingMready;�   5   7   L      +                        bitCounter    := 0;�   4   6   L      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   3   5   L      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   2   4   L      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   1   3   L      H                        index         := to_integer(unsigned(data2Map));�   0   2   L      \                     if bitCounter = 4 then                             --porque bit voy?   �   /   1   L      >                     bitCounter             := bitCounter + 2;�   .   0   L      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   -   /   L      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   ,   .   L      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   +   -   L      $               when waitingSvalid =>�   *   ,   L                  case state is�   )   +   L               else�   (   *   L      -            data2Map      <= (others => '0');�   '   )   L      -            m_axis_tdata  <= (others => '0');�   &   (   L      !            m_axis_tvalid <= '0';�   %   '   L      !            s_axis_tready <= '1';�   $   &   L      +            state         <= waitingSvalid;�   #   %   L               if rst = '0' then�   "   $   L            if rising_edge(clk) then�   !   #   L         begin�       "   L      1      variable index      :natural range 0 to 15;�      !   L      1      variable bitCounter :natural range 0 to 8 ;�          L      %   mapper_proc:process (clk) is --{{{�         L      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;�         L      2   signal state      : axiStates := waitingSvalid;�         L      4   type axiStates is (waitingSvalid, waitingMready);�         L      �   constant im_table   : real_im_array := (25 ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         L      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         L      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         L      *           rst           : in  STD_LOGIC);�         L      )           clk           : in  STD_LOGIC;�         L      )           s_axis_tready : out STD_LOGIC;�         L      )           s_axis_tlast  : in  STD_LOGIC;�         L      )           s_axis_tvalid : in  STD_LOGIC;�         L      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   	      L      )           m_axis_tready : in  STD_LOGIC;�      
   L      )           m_axis_tlast  : out STD_LOGIC;�      	   L      )           m_axis_tvalid : out STD_LOGIC;�         L      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         L          Port(  �                �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�                �   constant im_table   : real_im_array  := (25 ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^L�   d �   I   K   L      !   end process mapper_proc; --}}}�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L                     when others =>�   D   F   L                        end if;�   C   E   L                           end if;�   B   D   L      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   A   C   L      +                        bitCounter    := 0;�   @   B   L      -                        s_axis_tready <= '1';�   ?   A   L      �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   >   @   L                           else�   =   ?   L      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));�   <   >   L      a                     if bitCounter < 2 then                        --perfecto, porque bit voy?   �   ;   =   L      O                     bitCounter := bitCounter+1;                   --incremento�   :   <   L      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   9   ;   L      $               when waitingMready =>�   8   :   L                        end if;�   7   9   L                           end if;�   6   8   L      7                        state         <= waitingMready;�   5   7   L      +                        bitCounter    := 0;�   4   6   L      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   3   5   L      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   2   4   L      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   1   3   L      H                        index         := to_integer(unsigned(data2Map));�   0   2   L      \                     if bitCounter = 4 then                             --porque bit voy?   �   /   1   L      >                     bitCounter             := bitCounter + 2;�   .   0   L      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   -   /   L      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   ,   .   L      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   +   -   L      $               when waitingSvalid =>�   *   ,   L                  case state is�   )   +   L               else�   (   *   L      -            data2Map      <= (others => '0');�   '   )   L      -            m_axis_tdata  <= (others => '0');�   &   (   L      !            m_axis_tvalid <= '0';�   %   '   L      !            s_axis_tready <= '1';�   $   &   L      +            state         <= waitingSvalid;�   #   %   L               if rst = '0' then�   "   $   L            if rising_edge(clk) then�   !   #   L         begin�       "   L      1      variable index      :natural range 0 to 15;�      !   L      1      variable bitCounter :natural range 0 to 8 ;�          L      %   mapper_proc:process (clk) is --{{{�         L      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;�         L      2   signal state      : axiStates := waitingSvalid;�         L      4   type axiStates is (waitingSvalid, waitingMready);�         L      �   constant im_table   : real_im_array := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         L      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         L      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         L      *           rst           : in  STD_LOGIC);�         L      )           clk           : in  STD_LOGIC;�         L      )           s_axis_tready : out STD_LOGIC;�         L      )           s_axis_tlast  : in  STD_LOGIC;�         L      )           s_axis_tvalid : in  STD_LOGIC;�         L      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   	      L      )           m_axis_tready : in  STD_LOGIC;�      
   L      )           m_axis_tlast  : out STD_LOGIC;�      	   L      )           m_axis_tvalid : out STD_LOGIC;�         L      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         L          Port(  �                �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�                �   constant im_table   : real_im_array := (25 ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);5�_�  �  �          �   2   A    ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^N�     �   1   3   L      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^N�   e �       "   L      1      variable index      :natural range 0 to 15;5�_�  �  �          �   !   *    ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^P�     �       "   L    �   !   "   L    5�_�  �  �          �   "       ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^P�     �   !   #   M      1      variable index      :integer range 0 to 15;5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                               3          3       V   3    ^P�     �   /   1   M    �   0   1   M    5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          1          v       ^P�     �   0   2   N      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          1   &       v   &    ^P�   f �   0   2   N      ;                     test(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          1   &       v   &    ^P�     �   0   2   N      -                     test <= s_axis_tdata(1);5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          1   &       v   &    ^P�   g �   0   2   N      -                     test "= s_axis_tdata(1);5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          1   &       v   &    ^P�     �   0   2   N      -                     test := s_axis_tdata(1);5�_�  �  �          �   "       ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�     �   !   #   N      0      variable test      :integer range 0 to 15;5�_�  �  �  �      �   "   +    ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�     �   !   #   N      9      variable test      :std_logic_vector range 0 to 15;5�_�  �  �          �   "   +    ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�     �   !   #   N      +      variable test      :std_logic_vector 5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�   h �   0   2   N      .                     test( := s_axis_tdata(1);5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�   i �   0   2   N      0                     test(0) := s_axis_tdata(1);5�_�  �  �  �      �   1        ����                                                                                                                                                                                                                                                                                                                            /   5       0   5       V   5    ^Q     �   0   3   N    �   1   2   N    5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            1          2                 ^Q     �   0   2   P      7                     (bitCounter)   <= s_axis_tdata(0);�   0   3   P      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);   ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            1          2                 ^Q   j �   2   3          9                     test(bitCounter) := s_axis_tdata(1);5�_�  �  �  �      �   /        ����                                                                                                                                                                                                                                                                                                                            /          2          V       ^Q$   k �   L   N   O      !   end process mapper_proc; --}}}�   K   M   O            end if;�   J   L   O               end if;�   I   K   O                  end case;�   H   J   O                     when others =>�   G   I   O                        end if;�   F   H   O                           end if;�   E   G   O      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   D   F   O      +                        bitCounter    := 0;�   C   E   O      -                        s_axis_tready <= '1';�   B   D   O      �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   A   C   O                           else�   @   B   O      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));�   ?   A   O      a                     if bitCounter < 2 then                        --perfecto, porque bit voy?   �   >   @   O      O                     bitCounter := bitCounter+1;                   --incremento�   =   ?   O      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   <   >   O      $               when waitingMready =>�   ;   =   O                        end if;�   :   <   O                           end if;�   9   ;   O      7                        state         <= waitingMready;�   8   :   O      +                        bitCounter    := 0;�   7   9   O      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   6   8   O      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   5   7   O      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));�   4   6   O      H                        index         := to_integer(unsigned(data2Map));�   3   5   O      \                     if bitCounter = 4 then                             --porque bit voy?   �   2   4   O      >                     bitCounter             := bitCounter + 2;�   1   3   O      ?                     test(bitCounter+1)     <= s_axis_tdata(1);�   0   2   O      ?                     test(bitCounter)       <= s_axis_tdata(0);�   /   1   O      ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   .   0   O      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   -   /   O      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   ,   .   O      $               when waitingSvalid =>�   +   -   O                  case state is�   *   ,   O               else�   )   +   O      -            data2Map      <= (others => '0');�   (   *   O      -            m_axis_tdata  <= (others => '0');�   '   )   O      !            m_axis_tvalid <= '0';�   &   (   O      !            s_axis_tready <= '1';�   %   '   O      +            state         <= waitingSvalid;�   $   &   O               if rst = '0' then�   #   %   O            if rising_edge(clk) then�   "   $   O         begin�   !   #   O      8      variable test      :std_logic_vector (7 downto 0);�       "   O      1      variable index      :integer range 0 to 15;�      !   O      1      variable bitCounter :natural range 0 to 8 ;�          O      %   mapper_proc:process (clk) is --{{{�         O      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;�         O      2   signal state      : axiStates := waitingSvalid;�         O      4   type axiStates is (waitingSvalid, waitingMready);�         O      �   constant im_table   : real_im_array := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);�         O      �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);�         O      F   type real_im_array is array (0 to 15) of integer range -128 to 127;�         O      *           rst           : in  STD_LOGIC);�         O      )           clk           : in  STD_LOGIC;�         O      )           s_axis_tready : out STD_LOGIC;�         O      )           s_axis_tlast  : in  STD_LOGIC;�         O      )           s_axis_tvalid : in  STD_LOGIC;�         O      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   	      O      )           m_axis_tready : in  STD_LOGIC;�      
   O      )           m_axis_tlast  : out STD_LOGIC;�      	   O      )           m_axis_tvalid : out STD_LOGIC;�         O      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         O          Port(  �   .   0          ?                     data2Map(bitCounter)   <= s_axis_tdata(0);�   0   2          ;                     test(bitCounter)   <= s_axis_tdata(0);�   /   1          ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);�   1   3          ;                     test(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   1   ,    ����                                                                                                                                                                                                                                                                                                                            1   ,       2   ,          ,    ^Q3   l �   0   3   O      ?                     test(bitCounter)       <= s_axis_tdata(0);   ?                     test(bitCounter+1)     <= s_axis_tdata(1);5�_�  �  �          �   5   =    ����                                                                                                                                                                                                                                                                                                                            1   ,       2   ,          ,    ^Q<   m �   4   6   O      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   *   )    ����                                                                                                                                                                                                                                                                                                                            1   ,       2   ,          ,    ^QS     �   )   +   O    �   *   +   O    5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            2   ,       3   ,          ,    ^QT     �   *   ,   P      -            data2Map      <= (others => '0');5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            2   ,       3   ,          ,    ^QW   n �   *   ,   P      )            test      <= (others => '0');5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                            2   ,       3   ,          ,    ^Qe     �   6   8   P    �   7   8   P    5�_�  �  �          �   7   O    ����                                                                                                                                                                                                                                                                                                                            7   O       7   S       v   S    ^Qp   o �   6   8   Q      Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                            7   O       7   S       v   S    ^Q}   q �   6   7          Y                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(test),8));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       ^V�     �         P      7   signal data2Map   :std_logic_vector ( 7 downto 0 ) ;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                V       ^V�     �                9   variable data2Map   :std_logic_vector ( 7 downto 0 ) ;5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                            !           !           V        ^V�     �       "   N    �   !   "   N    �       !          8      variable test      :std_logic_vector (7 downto 0);5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            !           !   8       V        ^V�     �       "          9   variable data2Map   :std_logic_vector ( 7 downto 0 ) ;5�_�  �  �          �   *       ����                                                                                                                                                                                                                                                                                                                            !           !   8       V        ^V�     �   )   *          )            test      := (others => '0');5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            !           !   8       V        ^V�     �   (   *   N      -            data2Map      <= (others => '0');5�_�  �  �          �   0        ����                                                                                                                                                                                                                                                                                                                            0          1          V       ^V�     �   /   0          ?                     test(bitCounter)       := s_axis_tdata(0);   ?                     test(bitCounter+1)     := s_axis_tdata(1);5�_�  �  �          �   .   ,    ����                                                                                                                                                                                                                                                                                                                            /   ,       .   ,          ,    ^V�   r �   -   0   L      ?                     data2Map(bitCounter)   <= s_axis_tdata(0);   ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   .   ,    ����                                                                                                                                                                                                                                                                                                                            .   ,       /   ,          ,    ^V�   s �   -   0   L      ?                     data2Map(bitCounter)   '= s_axis_tdata(0);   ?                     data2Map(bitCounter+1) '= s_axis_tdata(1);5�_�  �              �   2   =    ����                                                                                                                                                                                                                                                                                                                            2   =       2   @       v   @    ^V�   t �   1   3   L      D                        index         := to_integer(unsigned(test));5�_�  �          �  �   0       ����                                                                                                                                                                                                                                                                                                                            2          0          V       ^Q!     �   /   3   O      ?kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk   ;kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk   ;kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                                                v       ^Q     �         N      1    data2Map   :std_logic_vector ( 7 downto 0 ) ;5�_�  �          �  �   "   +    ����                                                                                                                                                                                                                                                                                                                            "          "           v        ^P�     �   !   #   N      �      variable test      :std_logic_vector (7 downto 0(7 downto 0(7 downto 0(7 downto 0(7 downto 0(7 downto 0(7 downto 0(7 downto 0(7 downto 0range 0 to 15;5�_�  �  �      �  �           ����                                                                                                                                                                                                                                                                                                                                                  v        ^L�     �         L      �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �              �           ����                                                                                                                                                                                                                                                                                                                                                  v        ^L�     �         L      �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �  �      �  �   2       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�P     �   1   3   M      H                        index         := to_integer(unsigned(data2Map));5�_�  �  �          �   2   4    ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�U   [ �   1   3   M      R                        index         := to_integer("0101");--unsigned(data2Map));5�_�  �  �          �   2   <    ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�d   \ �   1   3   M      S                        index         := to_integer("0101"); --unsigned(data2Map));5�_�  �  �          �   2   4    ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�v     �   1   3   M      \                        index         := to_integer(unsigned("0101"); --unsigned(data2Map));5�_�  �  �          �   2   C    ����                                                                                                                                                                                                                                                                                                                            2   )       2   H       v   H    ^�z   ^ �   1   3   M      ]                        index         := to_integer(unsigned("0101")); --unsigned(data2Map));5�_�  �              �   2   )    ����                                                                                                                                                                                                                                                                                                                            2   )       2   H       v   H    ^��     �   1   3   M      N                        index         := lllllllllllllllllunsigned(data2Map));5�_�  �          �  �   2       ����                                                                                                                                                                                                                                                                                                                            )          %          V       ^�N     �   1   3        5�_�  �          �  �   ,       ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��     �   ,   -   L                           �   ,   .   M      '                     case bitCounter is   !                        when 0=> 5�_�  �          �  �   !   0    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^��   W �       "   K      3      variable index      :natural range 0 to 1500;5�_�  �  �      �  �   1   4    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�"     �   0   2   K      G                        index         := to_integer(nsigned(data2Map));5�_�  �              �   1   4    ����                                                                                                                                                                                                                                                                                                                            !   )       !   +       v   +    ^�"   U �   0   2   K      F                        index         := to_integer(signed(data2Map));5�_�  �      �  �  �   1   ,    ����                                                                                                                                                                                                                                                                                                                            :          D                 ^��     �   0   2   K      J                        index         := to_unsigned((unsigned(data2Map));5�_�  �          �  �   !   "    ����                                                                                                                                                                                                                                                                                                                            :          D                 ^�9   O �       "   K      5      variable index      :integer; -- range 0 to 15;5�_�  �  �      �  �   -       ����                                                                                                                                                                                                                                                                                                                            /          7                 ^��   H �   ,   .   K      A                     --data2Map(bitCounter)   <= s_axis_tdata(0);�   -   /   K      A                     --data2Map(bitCounter+1) <= s_axis_tdata(1);5�_�  �  �          �   /       ����                                                                                                                                                                                                                                                                                                                            /          7                 ^��   I �   .   0   K      @                     --bitCounter             := bitCounter + 2;�   /   8   K      ^                     --if bitCounter = 4 then                             --porque bit voy?      J                     --   index         := to_integer(unsigned(data2Map));   \                     --   m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   n                     --   s_axis_tready <= '0';                              --entonces yo tambien estoy listo   b                     --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada   -                     --   bitCounter    := 0;   9                     --   state         <= waitingMready;                        --end if;5�_�  �  �          �   -        ����                                                                                                                                                                                                                                                                                                                            0          8                 ^��     �   -   .   K    �   ,   -   K      !            m_axis_tvalid <= '0';5�_�  �  �          �   :       ����                                                                                                                                                                                                                                                                                                                            0          8                 ^��     �   :   ;   L    �   9   :   L      !            m_axis_tvalid <= '0';5�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                            0          8                 ^��     �   <   =   M    �   ;   <   M      !            m_axis_tvalid <= '0';5�_�  �              �   I       ����                                                                                                                                                                                                                                                                                                                            0          8                 ^��   J �   I   J   N    �   H   I   N      !            m_axis_tvalid <= '0';5�_�  �          �  �   #       ����                                                                                                                                                                                                                                                                                                                            #          G                 ^�2     �   "   $   J             00if rising_edge(clk) then�   #   H   J   $         00   if rst = '0' then   -      00      state         <= waitingSvalid;   #      00      s_axis_tready <= '1';   #      00      m_axis_tvalid <= '0';   /      00      m_axis_tdata  <= (others => '0');         00   else         00      case state is   &      00         when waitingSvalid =>   t      00            if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   A      00               data2Map(bitCounter)   <= s_axis_tdata(0);   A      00               data2Map(bitCounter+1) <= s_axis_tdata(1);   @      00               bitCounter             := bitCounter + 2;   ^      00               if bitCounter = 4 then                             --porque bit voy?      J      00                  index         := to_integer(unsigned(data2Map));   \      00                  m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   n      00                  s_axis_tready <= '0';                              --entonces yo tambien estoy listo   b      00                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada   -      00                  bitCounter    := 0;   9      00                  state         <= waitingMready;         00               end if;         00            end if;   &      00         when waitingMready =>   n      00            if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   Q      00               bitCounter := bitCounter+1;                   --incremento   c      00               if bitCounter < 2 then                        --perfecto, porque bit voy?      Z      00                  m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));         00               else   �      00                  m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   /      00                  s_axis_tready <= '1';   -      00                  bitCounter    := 0;         00                  state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato         00               end if;         00            end if;         00      end case;         00   end if;         00end if;5�_�  �      �  �  �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^9H     �         J      entity mapper is --{{{�         J      C           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0); --}}}5�_�  �          �  �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^8�     �         J      entity mapper is/*{{{*/�         J      end mapper;/*}}}*/5�_�  Q          S  R   0   @    ����                                                                                                                                                                                                                                                                                                                                                             ^/~     �   /   1   R      B                     bitCounter                 := bitCounter + 1;5�_�  ,          .  -   i   )    ����                                                                                                                                                                                                                                                                                                                            i   )       i   )       v   )    ^��     �   h   j   v      .                        m_axis_tdata  <= part;5�_�  #          %  $   ^        ����                                                                                                                                                                                                                                                                                                                            ^          c          V       ^�z     �   ]   d   u      Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Veeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   /eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �   �       �   �   5       ����                                                                                                                                                                                                                                                                                                                            5   "       5   1       v   1    ^��     �   4   6   L      z                     real_part := std_logic_vector(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �               �   5   "    ����                                                                                                                                                                                                                                                                                                                            5   "       5   1       v   1    ^��     �   4   6   L      q                     real_part := to_inge(to_signed(real_table(index),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �   �       �   �   2       ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^�t     �   1   3   I      8                     index := unsigned(s_axis_tdata),4);5�_�   �   �           �   2   4    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^�u     �   1   3   I      7                     index := unsigned(s_axis_tdata)4);5�_�   �   �           �   2   4    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^�u     �   1   3   I      6                     index := unsigned(s_axis_tdata));5�_�   �               �   2   4    ����                                                                                                                                                                                                                                                                                                                            2          2   (       v   (    ^�u   4 �   1   3   I      5                     index := unsigned(s_axis_tdata);5�_�   �           �   �   1   %    ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       v   %    ^��     �   0   2   F      y                     m_axis_tdata <= eTD_LOGIC_VECTOR(to_signed(real_table(1),8)); --to_integer(unsigned(s_axis_tdata)));5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                                v       ^�   # �         F      use IEEE.numeric_STDD.ALL;5�_�   �           �   �   1   <    ����                                                                                                                                                                                                                                                                                                                                                v       ^�x     �   0   2   F      a                     m_axis_tdata <= real_table(to_unsigned(ungiendhhhhhhhhhhhhhs_axis_tdata,4));5�_�   �           �   �   /       ����                                                                                                                                                                                                                                                                                                                               B          B          B    ^��     �   /   0   E    �   .   2   E      s                  if )s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   3                     )m_axis_tdata <= s_axis_tdata;                        5�_�   +           -   ,      2    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         A      8   signal mapper_table : mapper_array := (0=>x"12",1=>);5�_�                    )        ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^��     �   (   +   =      2eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   @eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5��