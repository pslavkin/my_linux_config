Vim�UnDo� � ��&��͝%R␊�xQ�D���}E��1O         N=1            g       g   g   g    ]�/s   
 _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(     �                 R//////////////////////////////////////////////////////////////////////////////////   // Module Name: lab1   R//////////////////////////////////////////////////////////////////////////////////    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(     �               module lab1(5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(     �               
enti lab1(5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(     �               entienti lab1(5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(%     �               entity lab1(5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�((     �               entity lab1 is(5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(3     �                  �             5�_�      	                 
    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(D     �                     port 5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(N     �                     generic N;5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(W     �                     N;5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(Z     �               	      N);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(]     �                     generic )5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(^     �                     generic *5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(m     �                     generic (5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(n     �                  generic (5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(n     �               	generic (5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(n     �               	generic (5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(n     �               	generic (5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(s     �                	generic (5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(v     �                      N5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(     �                     port ( 5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               
   port ( 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �                     input [3:0] swt,5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �                     swt input [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �                     swt in input [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �                     swt in [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �                      swt in std_loin [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               *      swt in std_logic_vectorin [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               )      swt in std_logic_vectorn [3:0] swt,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               (      swt in std_logic_vector [3:0] swt,5�_�                        "    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               '      swt in std_logic_vector[3:0] swt,5�_�      !                  "    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �               "      swt in std_logic_vector[3:0]5�_�       $           !      "    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�(�     �      	            �      	       5�_�   !   %   #       $          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)     �      	               led out std_;5�_�   $   &           %      #    ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)     �      	         %      led out std_logic_vector[3:0]_;5�_�   %   '           &   	       ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)     �      	                output [3:0] led5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)6     �               #      swt in std_logic_vector[3:0];5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                       ]�)8     �      	         $      swt in std_logic_vector [3:0];   $      led out std_logic_vector[3:0];5�_�   (   *           )           ����                                                                                                                                                                                                                                                                                                                                                          ]�)=     �               #      swt in std_logic_vector (30];�      	         $      swt in std_logic_vector (3:0];   $      led out std_logic_vector(3:0];5�_�   )   +           *      !    ����                                                                                                                                                                                                                                                                                                                               !          !          !    ]�)H     �      	         '      led out std_logic_vector(3 to 0];�               '      swt in std_logic_vector (3 to 0];5�_�   *   ,           +      )    ����                                                                                                                                                                                                                                                                                                                               )          )          )    ]�)O     �      	         +      swt in std_logic_vector (3 downto 0];   +      led out std_logic_vector(3 downto 0];5�_�   +   -           ,      )    ����                                                                                                                                                                                                                                                                                                                               )          )          )    ]�)Q     �      	         +      swt in std_logic_vector (3 downto 09;   +      led out std_logic_vector(3 downto 09;5�_�   ,   .           -      )    ����                                                                                                                                                                                                                                                                                                                               )          )          )    ]�)U     �      	         +      swt in std_logic_vector (3 downto 00;   +      led out std_logic_vector(3 downto 00;5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                               )          )          )    ]�)Z     �               +      swt in std_logic_vector (3 downto 0);5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                               )          )          )    ]�)[     �               ,      swt in  std_logic_vector (3 downto 0);5�_�   /   1           0           ����                                                                                                                                                                                                                                                                                                                                                V       ]�)\    �               $    assign led[3] = swt[2] & swt[3];�               $    assign led[2] = led[1] | led[3];�               %    assign led[1] = swt[1] & ~swt[2];�   
                assign led[0] = ~swt[0];�      
             );�      	         +      led out std_logic_vector(3 downto 0);�               +      swt in  std_logic_vector(3 downto 0);�               	   port (�                  );�                  N�                  generic (5�_�   0   2           1      	    ����                                                                                                                                                                                                                                                                                                                               	          	          	    ]�)e     �      	         .      led out std_logic_vector ( 3 downto 0 );�               .      swt in  std_logic_vector ( 3 downto 0 );5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                               	          	          	    ]�)q     �                  N5�_�   2   4           3   
        ����                                                                                                                                                                                                                                                                                                                               	          	          	    ]�)s     �   	             5�_�   3   5           4           ����                                                                                                                                                                                                                                                                                                                               	          	          	    ]�)x     �                5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                               	          	          	    ]�)�     �               end5�_�   5   7           6           ����                                                                                                                                                                                                                                                                                                                                         	       V       ]�)�     �                end   	endmodule5�_�   6   8           7           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)�     �                    assign led[0] = ~swt[0];   %    assign led[1] = swt[1] & ~swt[2];   $    assign led[2] = led[1] | led[3];   $    assign led[3] = swt[2] & swt[3];5�_�   7   9           8           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)�     �             �             5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �                    assign led[0] = ~swt[0];   %    assign led[1] = swt[1] & ~swt[2];   $    assign led[2] = led[1] | led[3];5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �               $    assign led[3] = swt[2] & swt[3];5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �                    led[3] = swt[2] & swt[3];5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �                    led[3] = swt[2] & swt[3];5�_�   <   >           =           ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �             �             5�_�   =   @           >          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �               end entity lab15�_�   >   A   ?       @          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �               end5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �               end entity lab5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �                �             5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               arquitecture 5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               arcuitecture 5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               archuitecture 5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               architecture 5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               architecture lab1_arq is 5�_�   G   I           H           ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �               !architecture lab1_arq of lab1 is 5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*     �                  �             5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*%     �               end entity lab15�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                V       ]�**    �               end architecture lab15�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*,     �               end architecture lab1_arq5�_�   L   N           M           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�*7     �               begin           end architecture lab1_arq;5�_�   M   O           N           ����                                                                                                                                                                                                                                                                                                                                                V       ]�*:     �   
            begin   end entity lab1;5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*>     �                  end entity lab1;5�_�   O   Q           P           ����                                                                                                                                                                                                                                                                                                                                                V       ]�*C    �                   end architecture lab1_arq;5�_�   P   R           Q           ����                                                                                                                                                                                                                                                                                                                                                V       ]�*r     �                 5�_�   Q   S           R      	    ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�     �               
use IEEE.;5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�     �               	use IEEE.5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�    �             5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�     �                5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�     �             �             5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                V       ]�*�     �             �             5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(3)<=0      led(3)<=0      led(3)<=05�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(2)<=0�                  led(2)<=0�                  led(2)<=05�_�   Y   [           Z          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(1)=swt(1)5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                   led(2)=1;5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(2)<=0      led(3)<=0      led(4)<=05�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(k)<=0      led(k)<=0      led(k)<=05�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(1)<=0�                  led(1)<=0�                  led(1)<=05�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(2)<=05�_�   _   a           `      	    ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(0)=swt(1)5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(0)<=swt(1)5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(1)<=05�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�     �                  led(2)<=15�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                       ]�*�    �                  led(3)<=05�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                                                       ]�-�    �                 5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                                                       ]�.T   	 �                 5�_�   f               g          ����                                                                                                                                                                                                                                                                                                                                                             ]�/r   
 �                  N=15�_�   >           @   ?          ����                                                                                                                                                                                                                                                                                                                                                V       ]�)�     �               end;   klu5�_�   !       "   $   #          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)     �      	         $      led out stdi   led out std_;_;5�_�   !           #   "          ����                                                                                                                                                                                                                                                                                                                                                  V        ]�)     �      	         #      led out std_   led out std_;;5��