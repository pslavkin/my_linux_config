Vim�UnDo� ��w�����Q\�F�[<�����?���̳��   =   2                     bitCounter := bitCounter + 8;   *   0                       ^$/�    _�                        1    ����                                                                                                                                                                                                                                                                                                                                                             ^$/�     �         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�                    )   -    ����                                                                                                                                                                                                                                                                                                                                                             ^$/�     �   (   *   =      R                     m_axis_tdata(bitCounter+7 downto bitCounter) <= s_axis_tdata;5�_�                     *   0    ����                                                                                                                                                                                                                                                                                                                                                             ^$/�    �   )   +   =      2                     bitCounter := bitCounter + 8;5��