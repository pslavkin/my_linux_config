Vim�UnDo� a6�쿅`;�H��.�wޭ�X|4x��yCg�2�3   L   2m_axis_config_tdata  <= "11111111"; --indirect FFT   I         H       H   H   H    ^))�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             ^&�<     �                +architecture Behavioral of slice_8from48 is�                end slice_8from48;�                entity slice_8from48 is5�_�                       1    ����                                                                                                                                                                                                                                                                                                                                                             ^&�H     �         G      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (47 downto 0);5�_�                    .   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   -   /   G      (                     bitCounter    := 0;5�_�                    .   (    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   -   /   G      *                     bitCounter    := 310;5�_�                    /   4    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   .   0   G      A                     m_axis_tdata  <= s_axis_tdata(37 downto 39);5�_�                    /   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   .   0   G      A                     m_axis_tdata  <= s_axis_tdata(30 downto 39);5�_�                    /   M    ����                                                                                                                                                                                                                                                                                                                                                             ^&�X     �   .   0   G      Q                     m_axis_tdata  <= (others=>'0') & s_axis_tdata(30 downto 39);5�_�      	              .   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   -   /   G      )                     bitCounter    := 31;5�_�      
           	   7   #    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   6   8   G      g                     if bitCounter < 16 then                             --perfecto, porque bit voy?   5�_�   	              
   7   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   6   8   G      g                     if bitCounter = 16 then                             --perfecto, porque bit voy?   5�_�   
                 9       ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   8   :   G                           else5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   8   :   G                           elsif�   9   :   G    5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   8   :   G      -                     elsifbitCounter = 1 then5�_�                    9   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   8   :   G      .                     elsif bitCounter = 1 then5�_�                    9   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   8   :   G    �   9   :   G    5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   8   :   H    �   9   :   H    5�_�                    :   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   9   ;   I      .                     elsif bitCounter = 2 then5�_�                   :   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   9   ;   I      .                     elsif bitCounter = r then5�_�                    ;   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   :   <   I      .                     elsif bitCounter = 2 then5�_�                    8   6    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�F     �   7   9   I      C                        m_axis_tdata  <= s_axis_tdata(14 downto 7);5�_�                    8   @    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�G     �   7   9   I      C                        m_axis_tdata  <= s_axis_tdata(23 downto 7);5�_�                    :   -    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�N     �   9   ;   I    �   :   ;   I    5�_�                    :   6    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�Q     �   9   ;   J      D                        m_axis_tdata  <= s_axis_tdata(23 downto 16);5�_�                    :   @    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�s     �   9   ;   J      D                        m_axis_tdata  <= s_axis_tdata(14 downto 16);5�_�                    :   @    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�t     �   9   ;   J      C                        m_axis_tdata  <= s_axis_tdata(14 downto 6);5�_�                    <   -    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�y     �   ;   =   J    �   <   =   J    5�_�                    <   6    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&�|     �   ;   =   K      C                        m_axis_tdata  <= s_axis_tdata(14 downto 8);5�_�                    <   ?    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   ;   =   K      B                        m_axis_tdata  <= s_axis_tdata(7 downto 8);5�_�                    :   )    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   9   ;   K      C                        m_axis_tdata  <= s_axis_tdata(14 downto 8);5�_�                     6   .    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   5   7   K      Q                     bitCounter := bitCounter+8;                     --incremento5�_�      !               =       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   <   >   K      .                     elsif bitCounter = 4 then5�_�       "           !   =       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   <   >   K                           els4 then5�_�   !   #           "   =       ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��    �   <   >   K                           elsen5�_�   "   $           #   /   &    ����                                                                                                                                                                                                                                                                                                                            /   &       /   0       v   0    ^&�     �   .   0   K      Q                     m_axis_tdata  <= (others=>'0') & s_axis_tdata(30 downto 24);5�_�   #   %           $   /   (    ����                                                                                                                                                                                                                                                                                                                            /   &       /   0       v   0    ^&�     �   .   0   K      G                     m_axis_tdata  <= "') & s_axis_tdata(30 downto 24);5�_�   $   &           %   /   )    ����                                                                                                                                                                                                                                                                                                                            /   &       /   0       v   0    ^&�     �   .   0   K      H                     m_axis_tdata  <= "'") & s_axis_tdata(30 downto 24);5�_�   %   '           &   /   '    ����                                                                                                                                                                                                                                                                                                                            /   &       /   0       v   0    ^&�    �   .   0   K      G                     m_axis_tdata  <= "'" & s_axis_tdata(30 downto 24);5�_�   &   (           '   :   )    ����                                                                                                                                                                                                                                                                                                                            :   )       :   2       v   2    ^&��     �   9   ;   K      S                        m_axis_tdata  <= (others=>'0') & s_axis_tdata(14 downto 8);5�_�   '   )           (   :   +    ����                                                                                                                                                                                                                                                                                                                            :   )       :   2       v   2    ^&��     �   9   ;   K      J                        m_axis_tdata  <= "0') & s_axis_tdata(14 downto 8);5�_�   (   *           )   :   ,    ����                                                                                                                                                                                                                                                                                                                            :   )       :   2       v   2    ^&��    �   9   ;   K      J                        m_axis_tdata  <= "0") & s_axis_tdata(14 downto 8);5�_�   )   +           *   :   +    ����                                                                                                                                                                                                                                                                                                                            :   )       :   2       v   2    ^&��    �   9   ;   K      I                        m_axis_tdata  <= "0" & s_axis_tdata(14 downto 8);5�_�   *   ,           +   :   +    ����                                                                                                                                                                                                                                                                                                                            :   )       :   2       v   2    ^&��    �   9   ;   K      J                        m_axis_tdata  <= "00" & s_axis_tdata(14 downto 8);5�_�   +   -           ,   F       ����                                                                                                                                                                                                                                                                                                                                                             ^&�9    �   F   H   K    5�_�   ,   .           -   /   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   .   0   L      G                     m_axis_tdata  <= "0" & s_axis_tdata(30 downto 24);5�_�   -   /           .   /   (    ����                                                                                                                                                                                                                                                                                                                                                             ^&��     �   .   0   L      G                     m_axis_tdata  <= '0" & s_axis_tdata(30 downto 24);5�_�   .   0           /   /   )    ����                                                                                                                                                                                                                                                                                                                                                             ^&��    �   .   0   L      G                     m_axis_tdata  <= '0' & s_axis_tdata(30 downto 24);5�_�   /   1           0   /   &    ����                                                                                                                                                                                                                                                                                                                                                             ^&�l     �   .   0   L      M                     m_axis_tdata  <= '0' & '0' & s_axis_tdata(30 downto 24);5�_�   0   2           1   /   (    ����                                                                                                                                                                                                                                                                                                                                                             ^&�n     �   .   0   L      O                     m_axis_tdata  <= x"'0' & '0' & s_axis_tdata(30 downto 24);5�_�   1   3           2   /   )    ����                                                                                                                                                                                                                                                                                                                                                             ^&�o     �   .   0   L      N                     m_axis_tdata  <= x"0' & '0' & s_axis_tdata(30 downto 24);5�_�   2   4           3   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�s     �   .   0   L      N                     m_axis_tdata  <= x"0" & '0' & s_axis_tdata(30 downto 24);5�_�   3   5           4   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�t     �   .   0   L      M                     m_axis_tdata  <= x"0"  '0' & s_axis_tdata(30 downto 24);5�_�   4   6           5   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�t     �   .   0   L      L                     m_axis_tdata  <= x"0" '0' & s_axis_tdata(30 downto 24);5�_�   5   7           6   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�u     �   .   0   L      K                     m_axis_tdata  <= x"0" 0' & s_axis_tdata(30 downto 24);5�_�   6   8           7   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�u     �   .   0   L      J                     m_axis_tdata  <= x"0" ' & s_axis_tdata(30 downto 24);5�_�   7   9           8   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^&�u     �   .   0   L      I                     m_axis_tdata  <= x"0"  & s_axis_tdata(30 downto 24);5�_�   8   :           9   :   )    ����                                                                                                                                                                                                                                                                                                                            :   )       :   0       v   0    ^&��     �   9   ;   L      N                        m_axis_tdata  <= "000000" & s_axis_tdata(14 downto 8);�   :   ;   L    5�_�   9   ;           :   :   0    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^&��     �   9   ;   L      M                        m_axis_tdata  <= x"0" &  & s_axis_tdata(14 downto 8);5�_�   :   <           ;   :   0    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^&��     �   9   ;   L      L                        m_axis_tdata  <= x"0" & & s_axis_tdata(14 downto 8);5�_�   ;   =           <   :   0    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^&��    �   9   ;   L      K                        m_axis_tdata  <= x"0" &  s_axis_tdata(14 downto 8);5�_�   <   >           =   :   )    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^&��     �   9   ;   L      J                        m_axis_tdata  <= x"0" & s_axis_tdata(14 downto 8);5�_�   =   ?           >   /   &    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^&�   
 �   .   0   L      H                     m_axis_tdata  <= x"0" & s_axis_tdata(30 downto 24);5�_�   >   @           ?   I        ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^'��     �   H   J   L      0m_axis_config_tdata  <= "00000000"; --direct FFT5�_�   ?   A           @   I   &    ����                                                                                                                                                                                                                                                                                                                            :   )       :   /       v   0    ^'��    �   H   J   L      0m_axis_config_tdata  <= "00000001"; --direct FFT5�_�   @   B           A   /   &    ����                                                                                                                                                                                                                                                                                                                            /   &       /   (       v   (    ^'�>     �   .   0   L      G                     m_axis_tdata  <= "0" & s_axis_tdata(30 downto 24);�   /   0   L    5�_�   A   C           B   /   2    ����                                                                                                                                                                                                                                                                                                                            /   &       /   1       v   (    ^'�?     �   .   0   L      P                     m_axis_tdata  <= s_axis_tdata & s_axis_tdata(30 downto 24);5�_�   B   D           C   :   )    ����                                                                                                                                                                                                                                                                                                                            :   )       :   +       v   +    ^'�P     �   9   ;   L      I                        m_axis_tdata  <= "0" & s_axis_tdata(14 downto 8);�   :   ;   L    5�_�   C   E           D   :   6    ����                                                                                                                                                                                                                                                                                                                            :   )       :   8       v   +    ^'�T     �   9   ;   L      V                        m_axis_tdata  <= s_axis_tdata(30) & s_axis_tdata(14 downto 8);5�_�   D   H           E   :   8    ����                                                                                                                                                                                                                                                                                                                            :   )       :   8       v   +    ^'�X    �   9   ;   L      V                        m_axis_tdata  <= s_axis_tdata(14l & s_axis_tdata(14 downto 8);5�_�   E       F       H   I        ����                                                                                                                                                                                                                                                                                                                            :   )       :   8       v   +    ^))�    �   H   J   L      2m_axis_config_tdata  <= "00000001"; --indirect FFT5�_�   E   G       H   F   I       ����                                                                                                                                                                                                                                                                                                                            :   )       :   8       v   +    ^'ڀ    �   H   J   L      2m_axis_config_tdata  <= "11111111"; --indirect FFT5�_�   F               G   I       ����                                                                                                                                                                                                                                                                                                                            :   )       :   8       v   +    ^'�!     �   H   J   L      2m_axis_config_tdata  <= "00000001"; --indirect FFT5�_�                    :   (    ����                                                                                                                                                                                                                                                                                                                            7          7   *       v   *    ^&��     �   9   ;   I      .                     elsif bitCounter = 4444en5��