Vim�UnDo� Kq��)���3�ʪhh�gQ{���+�廜Ӕ[   ?                 l       l   l   l    ^��    _�                            ����                                                                                                                                                                                                                                                                                                                                                             ^��     �         @      entity stretcher is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^�     �         @      end stretcher;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^�
    �         @      'architecture Behavioral of stretcher is5�_�                   /        ����                                                                                                                                                                                                                                                                                                                            0          6          V       ^��     �   .   6   @    �   /   0   @    5�_�                    8        ����                                                                                                                                                                                                                                                                                                                            8          9          V       ^��     �   7   8          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato   X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�                    2       ����                                                                                                                                                                                                                                                                                                                            8          8          V       ^��     �   1   2          T                        bitCounter      := bitCounter+1;                --incremento5�_�                    /       ����                                                                                                                                                                                                                                                                                                                            7          7          V       ^�     �   .   /          f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�                    1        ����                                                                                                                                                                                                                                                                                                                            1          3          V       ^�     �   0   1                               else   m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar5�_�                    /        ����                                                                                                                                                                                                                                                                                                                            /          0          V       ^�     �   /   1          X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   .   0          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    .        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�     �   =   ?   @         end process shift_reg;�   <   >   @            end if;�   ;   =   @               end if;�   :   <   @                  end case;�   9   ;   @                        end if;�   8   :   @      �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   7   9   @                        else�   6   8   @                           end if;�   5   7   @      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar�   4   6   @      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   3   5   @                           else�   2   4   @      T                        bitCounter      := bitCounter+1;                --incremento�   1   3   @      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   0   2   @      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   /   1   @      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   .   0   @      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   -   /   @      a                     s_axis_tready   <= '0';--el dato esta en la mesa, ya no quiero mas por ahora�   ,   .   @      $               when waitingMready =>�   +   -   @                        end if;�   *   ,   @      (                     bitCounter    := 0;�   )   +   @      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   (   *   @      i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo�   '   )   @      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   @      $               when waitingSvalid =>�   %   '   @                  case state is�   $   &   @               else�   #   %   @      -            m_axis_tdata  <= (others => '0');�   "   $   @      !            m_axis_tvalid <= '0';�   !   #   @      !            s_axis_tready <= '0';�       "   @      +            state         <= waitingSvalid;�      !   @               if rst = '0' then�          @            if rising_edge(clk) then�         @         begin�         @      0      variable bitCounter :integer range 0 to 8;�         @         shift_reg:process (clk) is�         @      ,   signal state:shiftState := waitingSvalid;�         @      5   type shiftState is (waitingSvalid, waitingMready);�         @      *           rst           : in  STD_LOGIC);�         @      )           clk           : in  STD_LOGIC;�         @      )           s_axis_tready : out STD_LOGIC;�         @      )           s_axis_tlast  : in  STD_LOGIC;�         @      )           s_axis_tvalid : in  STD_LOGIC;�         @      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         @      )           m_axis_tready : in  STD_LOGIC;�   
      @      )           m_axis_tlast  : out STD_LOGIC;�   	      @      )           m_axis_tvalid : out STD_LOGIC;�      
   @      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   @          Port(  �   -   /          }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   /   1          U                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   .   0          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    .   ,    ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�     �   -   /   @      a                     s_axis_tready   <= '0';--el dato esta en la mesa, ya no quiero mas por ahora5�_�      !               )       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�b     �   (   )          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�       "           !   -       ����                                                                                                                                                                                                                                                                                                                            -          /          V       ^�s     �   ,   -          z                     s_axis_tready   <= '0';                         --el dato esta en la mesa, ya no quiero mas por ahora5�_�   !   #           "   4        ����                                                                                                                                                                                                                                                                                                                            4           4           V        ^��     �   3   4          r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar5�_�   "   $           #   3       ����                                                                                                                                                                                                                                                                                                                            4           4           V        ^��     �   2   4   =    �   3   4   =    5�_�   #   %           $   3        ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   2   4   >      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar   m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�   $   &           %   4       ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   3   5   =    �   4   5   =    5�_�   %   '           &   4       ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   3   5          !            s_axis_tready <= '0';5�_�   &   )           '   4   *    ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   3   5   >      -                        s_axis_tready <= '0';5�_�   '   *   (       )   5       ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   4   6   >    �   5   6   >    5�_�   )   +           *   5       ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   4   6          �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   *   ,           +   5   0    ����                                                                                                                                                                                                                                                                                                                            5          5          V       ^��     �   4   6   ?      �                        state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   +   -           ,   7        ����                                                                                                                                                                                                                                                                                                                            7          8   5       V   5    ^�     �   6   7                            else   �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)5�_�   ,   .           -   0   %    ����                                                                                                                                                                                                                                                                                                                            7          7   5       V   5    ^��     �   /   1   =      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�   -   /           .   0   %    ����                                                                                                                                                                                                                                                                                                                            7          7   5       V   5    ^��     �   /   1   =      f                     if bitCounter < 7 then                             --perfecto, porque bit voy?   5�_�   .   0           /   1        ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �   0   1          T                        bitCounter      := bitCounter+1;                --incremento5�_�   /   1           0   0       ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �   /   1   <    �   0   1   <    5�_�   0   2           1   0       ����                                                                                                                                                                                                                                                                                                                            2   %       2   %       V   %    ^��     �   /   1   =      T                        bitCounter      := bitCounter+1;                --incremento5�_�   1   3           2   0       ����                                                                                                                                                                                                                                                                                                                            2   %       2   %       V   %    ^��     �   /   1   =      T                     q  bitCounter      := bitCounter+1;                --incremento5�_�   2   4           3   0       ����                                                                                                                                                                                                                                                                                                                            2   %       2   %       V   %    ^��     �   /   1   =      S                       bitCounter      := bitCounter+1;                --incremento5�_�   3   5           4   0       ����                                                                                                                                                                                                                                                                                                                            2   %       2   %       V   %    ^��     �   /   1   =      R                      bitCounter      := bitCounter+1;                --incremento5�_�   4   6           5   0        ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^��     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =                           end if;�   4   6   =      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   3   5   =      -                        s_axis_tready <= '1';�   2   4   =      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   1   3   =                           else�   0   2   =      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   /   1   =      <                     bitCounter := bitCounter+1;--incremento�   .   0   =      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   -   /   =      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   ,   .   =      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   +   -   =      $               when waitingMready =>�   *   ,   =                        end if;�   )   +   =      (                     bitCounter    := 0;�   (   *   =      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   '   )   =      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   =      $               when waitingSvalid =>�   %   '   =                  case state is�   $   &   =               else�   #   %   =      -            m_axis_tdata  <= (others => '0');�   "   $   =      !            m_axis_tvalid <= '0';�   !   #   =      !            s_axis_tready <= '0';�       "   =      +            state         <= waitingSvalid;�      !   =               if rst = '0' then�          =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         =      )           m_axis_tready : in  STD_LOGIC;�   
      =      )           m_axis_tlast  : out STD_LOGIC;�   	      =      )           m_axis_tvalid : out STD_LOGIC;�      
   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   =          Port(  �   /   1          Q                     bitCounter      := bitCounter+1;                --incremento5�_�   5   9           6   0   0    ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^��     �   /   1   =      <                     bitCounter := bitCounter+1;--incremento5�_�   6   :   7       9   -        ����                                                                                                                                                                                                                                                                                                                            -   #       -   #       V   #    ^�?     �   ,   -          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   9   ;           :   1       ����                                                                                                                                                                                                                                                                                                                            -   #       -   #       V   #    ^�A     �   0   2   <    �   1   2   <    5�_�   :   <           ;   1       ����                                                                                                                                                                                                                                                                                                                            -   #       -   #       V   #    ^�B     �   0   2          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   ;   =           <   -        ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^�y     �   ,   -          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   <   >           =   1       ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^�z     �   0   2   <    �   1   2   <    5�_�   =   ?           >   1       ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^�{     �   0   2          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   >   @           ?   0        ����                                                                                                                                                                                                                                                                                                                            0          1          V       ^��     �   /   0          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato   W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   ?   A           @   -       ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^��     �   ,   /   ;    �   -   .   ;    5�_�   @   B           A   -        ����                                                                                                                                                                                                                                                                                                                            -          .          V       ^��     �   -   /          W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   ,   .          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   A   C           B   1   #    ����                                                                                                                                                                                                                                                                                                                            -          .          V       ^��     �   0   2   =      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�   B   D           C   +        ����                                                                                                                                                                                                                                                                                                                            -   #       .   #       V   #    ^�i     �   *   -   =    �   +   ,   =    5�_�   C   E           D   +        ����                                                                                                                                                                                                                                                                                                                            +          ,          V       ^�j     �   +   -          Q                  m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   *   ,          n                  m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   D   F           E   /        ����                                                                                                                                                                                                                                                                                                                            /          0          V       ^�p     �   .   /          n                  m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato   Q                  m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   E   G           F   2       ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^�w     �   1   4   =    �   2   3   =    5�_�   F   H           G   2        ����                                                                                                                                                                                                                                                                                                                            2          3          V       ^�x     �   2   4          Q                  m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   1   3          n                  m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   G   I           H   1   #    ����                                                                                                                                                                                                                                                                                                                            2          3          V       ^��    �   0   2   ?      f                     if bitCounter = 8 then                             --perfecto, porque bit voy?   5�_�   H   J           I   *       ����                                                                                                                                                                                                                                                                                                                            2          3          V       ^��     �   )   +   ?    �   *   +   ?    5�_�   I   K           J   *       ����                                                                                                                                                                                                                                                                                                                            3          4          V       ^��     �   )   +          -                        s_axis_tready <= '1';5�_�   J   L           K   *   '    ����                                                                                                                                                                                                                                                                                                                            3          4          V       ^��     �   )   +   @      *                     s_axis_tready <= '1';5�_�   K   N           L   )        ����                                                                                                                                                                                                                                                                                                                            -   '       )   '       V   '    ^��     �   =   ?   @         end process shift_reg;�   <   >   @            end if;�   ;   =   @               end if;�   :   <   @                  end case;�   9   ;   @                        end if;�   8   :   @                           end if;�   7   9   @      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   6   8   @      -                        s_axis_tready <= '1';�   5   7   @      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   4   6   @                           else�   3   5   @      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   2   4   @      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   1   3   @      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   0   2   @      Q                     bitCounter := bitCounter+1;                     --incremento�   /   1   @      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   .   0   @      $               when waitingMready =>�   -   /   @                        end if;�   ,   .   @      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   +   -   @      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   *   ,   @      *                     bitCounter      := 0;�   )   +   @      ,                     s_axis_tready   <= '0';�   (   *   @      p                     state           <= waitingMready;--cambio de estado, y le doy un clk para que ponga el dato�   '   )   @      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   @      $               when waitingSvalid =>�   %   '   @                  case state is�   $   &   @               else�   #   %   @      -            m_axis_tdata  <= (others => '0');�   "   $   @      !            m_axis_tvalid <= '0';�   !   #   @      !            s_axis_tready <= '0';�       "   @      +            state         <= waitingSvalid;�      !   @               if rst = '0' then�          @            if rising_edge(clk) then�         @         begin�         @      0      variable bitCounter :integer range 0 to 8;�         @         shift_reg:process (clk) is�         @      ,   signal state:shiftState := waitingSvalid;�         @      5   type shiftState is (waitingSvalid, waitingMready);�         @      *           rst           : in  STD_LOGIC);�         @      )           clk           : in  STD_LOGIC;�         @      )           s_axis_tready : out STD_LOGIC;�         @      )           s_axis_tlast  : in  STD_LOGIC;�         @      )           s_axis_tvalid : in  STD_LOGIC;�         @      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         @      )           m_axis_tready : in  STD_LOGIC;�   
      @      )           m_axis_tlast  : out STD_LOGIC;�   	      @      )           m_axis_tvalid : out STD_LOGIC;�      
   @      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   @          Port(  �   (   *          �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   ,   .          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   +   -          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   *   ,          (                     bitCounter    := 0;�   )   +          *                     s_axis_tready <= '0';5�_�   L   O   M       N   )   6    ����                                                                                                                                                                                                                                                                                                                            -   '       )   '       V   '    ^��     �   (   *   @      p                     state           <= waitingMready;--cambio de estado, y le doy un clk para que ponga el dato5�_�   N   P           O   )        ����                                                                                                                                                                                                                                                                                                                            )   %       )   %       V   %    ^��     �   (   )                               state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato5�_�   O   Q           P   -       ����                                                                                                                                                                                                                                                                                                                            )   %       )   %       V   %    ^      �   ,   .   ?    �   -   .   ?    5�_�   P   R           Q   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^ 
     �   +   ,          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   Q   S           R   +       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^     �   *   ,   ?    �   +   ,   ?    5�_�   R   T           S   3       ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^ Z    �   2   3          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   S   U           T   "       ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^'    �   !   #   ?      !            s_axis_tready <= '0';5�_�   T   V           U   +   <    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   *   ,   ?    �   +   ,   ?    5�_�   U   W           V   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   +   -   @    �   ,   -   @    5�_�   V   X           W   -   "    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   ,   .   A      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   W   Y           X   -   ?    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   ,   .   A      T                     m_axis_tdata(1) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   X   Z           Y   +       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   *   ,   A      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   Y   [           Z   3   -    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   2   4   A    �   3   4   A    5�_�   Z   \           [   3       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   2   4   B      Q                     bitCounter := bitCounter+1;                     --incremento5�_�   [   ]           \   4   .    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   3   5   B      Q                     bitCounter := bitCounter+1;                     --incremento5�_�   \   ^           ]   6   .    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   5   7   B    �   6   7   B    5�_�   ]   _           ^   7   %    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   6   8   C      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   ^   `           _   7   B    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   6   8   C      W                        m_axis_tdata(1) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   _   a           `   6   B    ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   5   7   C    �   6   7   C    5�_�   `   b           a   6       ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   5   7   D      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   a   c           b   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   +   ,          T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   b   d           c   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   +   ,          V                     m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�   c   e           d   +       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   *   ,   B      V                     --m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   d   f           e   +       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   *   ,   B      U                     -m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   e   g           f   2       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   1   2          Q                     bitCounter := bitCounter+2;                     --incremento5�_�   f   h           g   1       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   0   2   A      S                     --bitCounter := bitCounter+1;                     --incremento5�_�   g   j           h   1       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   0   2   A      R                     -bitCounter := bitCounter+1;                     --incremento5�_�   h   k   i       j   3       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   2   4   A      Y                        --m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   j   l           k   3       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   2   4   A      X                        -m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�   k               l   4        ����                                                                                                                                                                                                                                                                                                                            4          5          V       ^��    �   3   4          W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato   Y                        m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�   h           j   i   3       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   2   4        5�_�   L           N   M   )   6    ����                                                                                                                                                                                                                                                                                                                            .   '       )   '       V   '    ^��     �   )   *   @       5�_�   6   8       9   7   1   #    ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^�     �   0   2   =      f                     if bitCounter = 8 then                             --perfecto, porque bit voy?   5�_�   7               8   2       ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^�     �   1   3        5�_�   '           )   (   5       ����                                                                                                                                                                                                                                                                                                                            3          3          V       ^��     �   5   6   >    �   5   6   >      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�                    .   ,    ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�     �   -   /   @      �                     s_axis_tready   <= '0';                         hhhhhhhhhhhhhhhhhhhhhhhhhhhh--el dato esta en la mesa, ya no quiero mas por ahora5�_�                   /       ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^��     �   /   0   @    �   .   /   @      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    /       ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^��     �   .   0          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    /   #    ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^��     �   .   0   A      p                     m_axis_tvalid  <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    /   #    ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^��     �   .   0   A      o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�      	              .       ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^�>     �   -   /        5�_�      
           	   1       ����                                                                                                                                                                                                                                                                                                                            '           ,           V        ^�?     �   1   2   @    �   0   1   @      }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�   	              
   1       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^�A     �   0   2          �                        s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�   
                 1        ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^�B     �   0   2        5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^�F     �   0   1   @    �   /   0   @      �                        s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^�H     �   -   /        5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^��     �   )   *   @    �   (   )   @      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            *   '       )   '       V   '    ^��     �   (   *          U                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�                    )        ����                                                                                                                                                                                                                                                                                                                            )          ,          V       ^��     �   )   +          k                     s_axis_tready   <= '1';                              --entonces yo tambien estoy listo�   (   *          P                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);--pongo el dato�      	   A          Port(  �      
   A      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   	      A      )           m_axis_tvalid : out STD_LOGIC;�   
      A      )           m_axis_tlast  : out STD_LOGIC;�         A      )           m_axis_tready : in  STD_LOGIC;�         A      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         A      )           s_axis_tvalid : in  STD_LOGIC;�         A      )           s_axis_tlast  : in  STD_LOGIC;�         A      )           s_axis_tready : out STD_LOGIC;�         A      )           clk           : in  STD_LOGIC;�         A      *           rst           : in  STD_LOGIC);�         A      5   type shiftState is (waitingSvalid, waitingMready);�         A      ,   signal state:shiftState := waitingSvalid;�         A         shift_reg:process (clk) is�         A      0      variable bitCounter :integer range 0 to 8;�         A         begin�          A            if rising_edge(clk) then�      !   A               if rst = '0' then�       "   A      +            state         <= waitingSvalid;�   !   #   A      !            s_axis_tready <= '0';�   "   $   A      !            m_axis_tvalid <= '0';�   #   %   A      -            m_axis_tdata  <= (others => '0');�   $   &   A               else�   %   '   A                  case state is�   &   (   A      $               when waitingSvalid =>�   '   )   A      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   (   *   A      P                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);--pongo el dato�   )   +   A      k                     s_axis_tready   <= '1';                              --entonces yo tambien estoy listo�   *   ,   A      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   +   -   A      (                     bitCounter    := 0;�   ,   .   A                        end if;�   -   /   A      $               when waitingMready =>�   .   0   A      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   /   1   A      �                        s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   0   2   A      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   1   3   A      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   2   4   A      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   3   5   A      T                        bitCounter      := bitCounter+1;                --incremento�   4   6   A                           else�   5   7   A      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   6   8   A      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar�   7   9   A                           end if;�   8   :   A                        else�   9   ;   A      �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   :   <   A                        end if;�   ;   =   A                  end case;�   <   >   A               end if;�   =   ?   A            end if;�   >   @   A         end process shift_reg;5�_�                    )        ����                                                                                                                                                                                                                                                                                                                            )          ,          V       ^��     �   )   +          k                     s_axis_tready   <= '1';                              --entonces yo tambien estoy listo�   *   ,          �                     state           <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   +   -          *                     bitCounter      := 0;�   (   *          P                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);--pongo el dato�      	   A          Port(  �      
   A      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   	      A      )           m_axis_tvalid : out STD_LOGIC;�   
      A      )           m_axis_tlast  : out STD_LOGIC;�         A      )           m_axis_tready : in  STD_LOGIC;�         A      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         A      )           s_axis_tvalid : in  STD_LOGIC;�         A      )           s_axis_tlast  : in  STD_LOGIC;�         A      )           s_axis_tready : out STD_LOGIC;�         A      )           clk           : in  STD_LOGIC;�         A      *           rst           : in  STD_LOGIC);�         A      5   type shiftState is (waitingSvalid, waitingMready);�         A      ,   signal state:shiftState := waitingSvalid;�         A         shift_reg:process (clk) is�         A      0      variable bitCounter :integer range 0 to 8;�         A         begin�          A            if rising_edge(clk) then�      !   A               if rst = '0' then�       "   A      +            state         <= waitingSvalid;�   !   #   A      !            s_axis_tready <= '0';�   "   $   A      !            m_axis_tvalid <= '0';�   #   %   A      -            m_axis_tdata  <= (others => '0');�   $   &   A               else�   %   '   A                  case state is�   &   (   A      $               when waitingSvalid =>�   '   )   A      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   (   *   A      P                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);--pongo el dato�   )   +   A      k                     s_axis_tready   <= '1';                              --entonces yo tambien estoy listo�   *   ,   A      �                     state           <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato�   +   -   A      *                     bitCounter      := 0;�   ,   .   A                        end if;�   -   /   A      $               when waitingMready =>�   .   0   A      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   /   1   A      �                        s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   0   2   A      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   1   3   A      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   2   4   A      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   3   5   A      T                        bitCounter      := bitCounter+1;                --incremento�   4   6   A                           else�   5   7   A      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   6   8   A      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar�   7   9   A                           end if;�   8   :   A                        else�   9   ;   A      �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   :   <   A                        end if;�   ;   =   A                  end case;�   <   >   A               end if;�   =   ?   A            end if;�   >   @   A         end process shift_reg;5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^��     �   *   +   A    �   )   *   A      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^��     �   )   +          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    1        ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^��     �   0   2        5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^��     �   0   1   A    �   /   0   A      �                        s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�                     0       ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^��     �   /   1          z                  s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5��