Vim�UnDo� uĩ�p�*��S�u߀[��eہ_��+�{*/   =       aaa: component lab1   3                           ]��U    _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ]��%     �         %    �         %    5�_�                           ����                                                                                                                                                                                                                                                                                                                                       $           V        ]��'     �         ,        component design_1 is5�_�                            ����                                                                                                                                                                                                                                                                                                                                       $           V        ]��?     �      (   %    �         %    �                  component lab1 is     port (       reset_rtl : in STD_LOGIC;       sys_clock : in STD_LOGIC;       clk_out1 : out STD_LOGIC     );     end component design_1;5�_�                    (        ����                                                                                                                                                                                                                                                                                                                                       '          V        ]��M     �   '   )   /    �   (   )   /    5�_�                    (       ����                                                                                                                                                                                                                                                                                                                                       '          V        ]��O    �   '   )   0         end component;5�_�                    0        ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]��i     �   /   :   0    �   0            5�_�                    0       ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]��t     �   /   1   :         aaa:lab15�_�      	              5       ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]���     �   4   6   :                     clk=>clk_tb,5�_�      
           	   6       ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]���     �   5   7   :                     rst=>rst_tb,5�_�   	              
   6       ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]���     �   5   7   :                     rst=>'0',5�_�   
                 6       ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]���     �   5   7   :                     rst=>reset_rtl',5�_�                            ����                                                                                                                                                                                                                                                                                                                            *          /          V       ]��     �         :    �         :    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]��!     �         <      /      swt: in  std_logic_vector ( 2 downto 0 );   .      led: out std_logic_vector ( 3 downto 0 )5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]��$     �         <      ,    led: out std_logic_vector ( 3 downto 0 )�         <      -    swt: in  std_logic_vector ( 2 downto 0 );5�_�                      0    ����                                                                                                                                                                                                                                                                                                                                                       ]��+     �         <      0    led_rtl: out std_logic_vector ( 3 downto 0 )5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            9          :                 ]��5    �   8   :   <                     swt=>swt_,�   8   ;   <                     swt=>swt_tb,                  led=>led_tb5�_�                    .        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ]��I     �   :   <   <                  );�   9   ;   <                     led=>led_rtl�   8   :   <                     swt=>swt_rtl,�   7   9   <                     rst=>reset_rtl,�   6   8   <                     clk=>clk_1,�   5   7   <         port map (�   4   6   <                     )�   3   5   <                        N => 4�   2   4   <         generic map (�   1   3   <          aaa: component lab1�   0   2   <          );�   /   1   <            sys_clock => sys_clock�   .   0   <            reset_rtl => reset_rtl,�   -   /   <            clk_out1  => clk_out1,�   ,   .   <           port map (�   )   +   <         end component lab1;�   (   *   <          );�   '   )   <      .      led: out std_logic_vector ( 3 downto 0 )�   &   (   <      /      swt: in  std_logic_vector ( 2 downto 0 );�   %   '   <            clk: in  std_logic;�   $   &   <            rst: in  std_logic;�   #   %   <      	   port (�   "   $   <         );�   !   #   <                    N: natural :=1�       "   <         generic (�      !   <         component lab1 is�          <        end component design_1;�         <        );�         <          clk_out1 : out STD_LOGIC�         <          sys_clock : in STD_LOGIC;�         <          reset_rtl : in STD_LOGIC;�         <        port (�         <        component design_1 is�         <        );�         <          sys_clock : in STD_LOGIC�         <          reset_rtl : in STD_LOGIC;�         <          clk_out1 : out STD_LOGIC;�         <      1    led_rtl: out std_logic_vector ( 3 downto 0 );�         <      1    swt_rtl: in  std_logic_vector ( 2 downto 0 );�         <        port (�      	   <       --Purpose     : IP block netlist�         <       --Design      : design_1_wrapper�         <      3--Command     : generate_target design_1_wrapper.bd�         <      ,--Host        : work1 running 64-bit unknown�         <      (--Date        : Mon Nov  4 01:14:20 2019�   /   1                sys_clock => sys_clock�   .   0                reset_rtl => reset_rtl,�   -   /                clk_out1 => clk_out1,5�_�                    1        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ]��O    �   1   3   <    5�_�                     3        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ]��T    �   2   4   =          aaa: component lab15�_�                       /    ����                                                                                                                                                                                                                                                                                                                                                       ]��)     �         <      0    led_rtl: out std_logic_vector ( 3 downto 0 ;5��