Vim�UnDo� 5�v	%�K!1�l`�x��k�q_F�=.����c   Q   "               axi+s_tready<= '0';   =                      ^(�   4 _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ^|$     �                 R----------------------------------------------------------------------------------   -- Company:    -- Engineer:    --    &-- Create Date: 01/01/2020 07:49:01 AM   -- Design Name:    )-- Module Name: paralell2axi - Behavioral   -- Project Name:    -- Target Devices:    -- Tool Versions:    -- Description:    --    -- Dependencies:    --    -- Revision:   -- Revision 0.01 - File Created   -- Additional Comments:   --    R----------------------------------------------------------------------------------        5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ^|&     �                7-- Uncomment the following library declaration if using   6-- arithmetic functions with Signed or Unsigned values   --use IEEE.NUMERIC_STD.ALL;       ?-- Uncomment the following library declaration if instantiating   &-- any Xilinx leaf cells in this code.   --library UNISIM;   --use UNISIM.VComponents.all;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ^|,     �               #           m_last : out STD_LOGIC);�               "           m_ready : in STD_LOGIC;�   
            #           m_valid : out STD_LOGIC;�   	            !           s_last : in STD_LOGIC;�      
         #           s_ready : out STD_LOGIC;�      	         "           s_valid : in STD_LOGIC;�               4           emi : out STD_LOGIC_VECTOR (15 downto 0);�               3    Port ( emo : in STD_LOGIC_VECTOR (15 downto 0);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^|.     �               M    Port           ( emo :                in  STD_LOGIC_VECTOR (15 downto 0);5�_�                          ����                                                                                                                                                                                                                                                                                                                                                  V        ^|4     �               E    Port   ( emo :                in  STD_LOGIC_VECTOR (15 downto 0);5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                  V        ^|5     �               B    Port( emo :                in  STD_LOGIC_VECTOR (15 downto 0);5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  V        ^|9     �               C    Port(  emo :                in  STD_LOGIC_VECTOR (15 downto 0);5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^|;     �               $           m_last  : out STD_LOGIC);�               #           m_ready : in  STD_LOGIC;�               #           m_valid : out STD_LOGIC;�   
            #           s_last  : in  STD_LOGIC;�   	            #           s_ready : out STD_LOGIC;�      
         #           s_valid : in  STD_LOGIC;�      	         B           emi     : out STD_LOGIC_VECTOR (15 downto           0);�               C           emo :                in  STD_LOGIC_VECTOR (15 downto 0);�                   Port(  5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^|O     �               8           emo     : in  STD_LOGIC_VECTOR (15 downto 0);5�_�   
                        ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^|Q     �               9           emio     : in  STD_LOGIC_VECTOR (15 downto 0);5�_�                           ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^|R     �                8           emi     : out STD_LOGIC_VECTOR (15 downto 0);5�_�                            ����                                                                                                                                                                                                                                                                                                                                      
          V       ^|`     �                #           s_valid : in  STD_LOGIC;   #           s_ready : out STD_LOGIC;   #           s_last  : in  STD_LOGIC;5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                V       ^|c     �   	          �   
          5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|d     �   
            $           m_last  : out STD_LOGIC);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|f     �   
            #           m_clk  : out STD_LOGIC);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|l     �      	       �      	       5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	          V       ^|m     �      	         #           m_valid : out STD_LOGIC;5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	          V       ^|q     �      	         "           m_data : out STD_LOGIC;5�_�                       "    ����                                                                                                                                                                                                                                                                                                                            	          	          V       ^|u     �      	         #           m_data  : out STD_LOGIC;5�_�                            ����                                                                                                                                                                                                                                                                                                                            	          	          V       ^|�     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                            	          	          V       ^|�     �                  m_valid <= 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                  m_valid <=  emio (�                  m_data <= emio(7 downto 0);�               $           m_clk   : out STD_LOGIC);�   
            $           m_last  : out STD_LOGIC);�   	            #           m_ready : in  STD_LOGIC;�      
         #           m_valid : out STD_LOGIC;�      	         7           m_data  : out STD_LOGIC_VECTOR (7 downto 0);�               8           emio    : in  STD_LOGIC_VECTOR (15 downto 0);�                   Port(  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                  m_valid <= emio (5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                  m_valid <= emio(5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �   
             $           m_last  : out STD_LOGIC);5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �   	          �   
          5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                $           m_clk   : out STD_LOGIC);5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �   
          �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �             �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �             �             5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �             �             5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                  m_valid <= emio(8);5�_�   !   #           "      
    ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �                  m_last <= emio(8);5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �               8           emio    : in  STD_LOGIC_VECTOR (15 downto 0);5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                V       ^|�     �               <           emio    : inoout  STD_LOGIC_VECTOR (15 downto 0);5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                V       ^}     �                  m_valid <= emio(8);�                  m_valid <= emio(8);�                  m_last  <= emio(8);�                  m_valid <= emio(8);�                  m_data  <= emio(7 downto 0);�               #           m_ready : in  STD_LOGIC;�   
            $           m_clk   : out STD_LOGIC);�   	            $           m_last  : out STD_LOGIC);�      
         #           m_valid : out STD_LOGIC;�      	         7           m_data  : out STD_LOGIC_VECTOR (7 downto 0);�               ;           emio    : inout  STD_LOGIC_VECTOR (15 downto 0);�                   Port(  5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                V       ^},     �                  m_last  <= emio(8);5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                V       ^}1     �                  m_valid <= emio(8);5�_�   '   )           (      	    ����                                                                                                                                                                                                                                                                                                                                                V       ^}3     �                  m_clk <= emio(8);5�_�   (   +           )          ����                                                                                                                                                                                                                                                                                                                                                V       ^}5     �                  m_clk   <= emio(8);5�_�   )   ,   *       +          ����                                                                                                                                                                                                                                                                                                                                                V       ^};     �                  m_valid <= emio(8);5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                V       ^}D     �                  m_ready <= emio(8);5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                V       ^}P     �               "   emio(10) <= m_ready <= emio(8);5�_�   -   /           .           ����                                                                                                                                                                                                                                                                                                                                                V       ^}R     �                  emio(10) <= m_ready;�                  m_clk    <= emio(10);�                  m_last   <= emio(9);�                  m_valid <= emio(8);�                  m_data  <= emio(7 downto 0);�               %           m_ready : in    STD_LOGIC;�   
            &           m_clk   : out   STD_LOGIC);�   	            &           m_last  : out   STD_LOGIC);�      
         %           m_valid : out   STD_LOGIC;�      	         :           m_data  : out   STD_LOGIC_VECTOR (7  downto 0);�               :           emio    : inout STD_LOGIC_VECTOR (15 downto 0);�                   Port(  �                   emio(10) <= m_ready;�                   m_clk   <= emio(10);�                   m_last  <= emio(9);5�_�   .   0           /           ����                                                                                                                                                                                                                                                                                                                                                V       ^}X    �                 5�_�   /   1           0   
   $    ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^~�     �   	            &           m_last  : out   STD_LOGIC);   &           m_clk   : out   STD_LOGIC);5�_�   0   4           1      $    ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^~�    �               %           m_ready : in    STD_LOGIC;5�_�   1   5   2       4          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �               :           emio    : inout STD_LOGIC_VECTOR (15 downto 0);5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �               9           emio    : inut STD_LOGIC_VECTOR (15 downto 0);5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �               8           emio    : int STD_LOGIC_VECTOR (15 downto 0);5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �               7           emio    : in STD_LOGIC_VECTOR (15 downto 0);5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �               6           emi    : in STD_LOGIC_VECTOR (15 downto 0);5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^��     �             �             5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                               $          $          $    ^��     �      	         7           emi     : in STD_LOGIC_VECTOR (15 downto 0);5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                               $          $          $    ^��     �      	         7           emo     : in STD_LOGIC_VECTOR (15 downto 0);5�_�   ;   =           <           ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                  emio(10) <= m_ready;�                  m_clk    <= emio(10);�                  m_last   <= emio(9);�                  m_valid  <= emio(8);�                   m_data   <= emio(7 downto 0);�               &           m_ready : in    STD_LOGIC);�               %           m_clk   : out   STD_LOGIC;�   
            %           m_last  : out   STD_LOGIC;�   	            %           m_valid : out   STD_LOGIC;�      
         :           m_data  : out   STD_LOGIC_VECTOR (7  downto 0);�      	         8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�               7           emi     : in STD_LOGIC_VECTOR (15 downto 0);�                   Port(  5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                   m_data   <= emio(7 downto 0);5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                  m_valid  <= emio(8);5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                  m_last   <= emio(9);5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                  m_clk    <= emio(10);5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �                  emio(10) <= m_ready;5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                V       ^��    �                  emo(10) <= m_ready;5�_�   B   D           C           ����                                                                                                                                                                                                                                                                                                                            	                    V       ^��     �             �             5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                            	                    V       ^��     �             5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                       ^��     �               8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);   #           m_valid : out STD_LOGIC;   #           m_last  : out STD_LOGIC;   #           m_clk   : out STD_LOGIC;   $           m_ready : in  STD_LOGIC);5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                                       ^��     �               8           s_data  : out STD_LOGIC_VECTOR (7  downto 0);5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                       ^��     �               #           s_valid : out STD_LOGIC;5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               #           s_last  : out STD_LOGIC;5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                       ^�A     �               #           m_clk   : out STD_LOGIC;5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                                                       ^�B     �               "           _clk   : out STD_LOGIC;5�_�   J   L           K           ����                                                                                                                                                                                                                                                                                                                                                V       ^�C     �                !           clk   : out STD_LOGIC;5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                V       ^�E     �             �             5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                                                V       ^�F     �                #           s_clk   : out STD_LOGIC;5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                V       ^�H     �               $           s_ready : in  STD_LOGIC);5�_�   N   P           O           ����                                                                                                                                                                                                                                                                                                                                                V       ^�P     �                  emo(10)  <= m_ready;�                  m_clk    <= emi(10);�                  m_last   <= emi(9);�                  m_valid  <= emi(8);�                  m_data   <= emi(7 downto 0);�               #           clk     : out STD_LOGIC;�               $           s_ready : out STD_LOGIC);�               #           s_last  : in  STD_LOGIC;�               "           s_valid : in STD_LOGIC;�               8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�               $           m_ready : in  STD_LOGIC);�   
            #           m_last  : out STD_LOGIC;�   	            #           m_valid : out STD_LOGIC;�      
         8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	         8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�               8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�                   Port(  �                !           clk   : out STD_LOGIC;�                %           s_ready : out  STD_LOGIC);�                "           s_last  : in STD_LOGIC;�                7           s_data  : in STD_LOGIC_VECTOR (7  downto 0);�   
             #           m_last  : out STD_LOGIC;�   	             #           m_valid : out STD_LOGIC;�                $           m_ready : in  STD_LOGIC);5�_�   O   Q           P           ����                                                                                                                                                                                                                                                                                                                                                V       ^�T     �             5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                V       ^�U     �                  m_clk    <= emi(10);5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                                V       ^�U     �                  _clk    <= emi(10);5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                                                V       ^�V     �                   clk    <= emi(10);5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                V       ^�W     �             �               5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                                                V       ^�\     �      !       �             5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                                                V       ^�^     �       "   "    5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                V       ^�a     �         #         m_data   <= emi(7 downto 0);5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                                                V       ^�d     �         #         s_data   <= emi(7 downto 0);5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                V       ^�i     �         #      &   emo <= s_data   <= emi(7 downto 0);5�_�   Y   [           Z          ����                                                                                                                                                                                                                                                                                                                                                V       ^�q     �         #      2   emo(7 downto 0) <= s_data   <= emi(7 downto 0);5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                                V       ^�t     �         #         emo(7 downto 0) <= s_data;5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         #         m_valid  <= emi(8);5�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         #         emo(12m_valid  <= emi(8);5�_�   ]   _           ^      	    ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         #         emo(11m_valid  <= emi(8);5�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         #      !   emo(11) <= m_valid  <= emi(8);5�_�   _   a           `          ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �         #      !   emo(11) <= s_valid  <= emi(8);5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �          #         m_last   <= emi(9);�          #    5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �          #         emo(11) m_last   <= emi(9);5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �          #      !   emo(11) <= m_last   <= emi(9);5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �          #      !   emo(11) <= s_last   <= emi(9);5�_�   d   g           e          ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �          #      !   emo(12) <= s_last   <= emi(9);5�_�   e   h   f       g           ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �      !   #         emo(10)  <= m_ready;5�_�   g   i           h           ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �      !   #      "   s_ready <= emo(10)  <= m_ready;5�_�   h   j           i           ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �      !   #      "   s_ready <= emi(10)  <= m_ready;5�_�   i   k           j           ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �      !   #      "   s_ready <= emi(13)  <= m_ready;5�_�   j   l           k   "       ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �   !   #   #         clk    <= emi(10);5�_�   k   m           l   "       ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �   !   #   #         clk    <= emi(15);5�_�   l   n           m           ����                                                                                                                                                                                                                                                                                                                            "                    V       ^��     �   !   #   #         clk     <=     emi(14);�      !   #         s_ready <=     emi(13);�          #         emo(12) <=     s_last;�         #         emo(11) <=     s_valid;�         #      1   emo(7   downto 0)    <=     s_data(7 downto 0;�         #         emo(10) <=     m_ready;�         #         m_last  <=     emi(9);�         #         m_valid <=     emi(8);�         #      "   m_data  <=     emi(7 downto 0);�         #      #           clk     : out STD_LOGIC;�         #      $           s_ready : out STD_LOGIC);�         #      #           s_last  : in  STD_LOGIC;�         #      #           s_valid : in  STD_LOGIC;�         #      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         #      $           m_ready : in  STD_LOGIC);�   
      #      #           m_last  : out STD_LOGIC;�   	      #      #           m_valid : out STD_LOGIC;�      
   #      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   #      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         #      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         #          Port(  �                (   emo(7 downto 0) <= s_data(7 downto 0;�                   m_data   <= emi(7 downto 0);�                   emo(11) <= s_valid;�                   m_valid  <= emi(8);�                    emo(12) <= s_last;�      !             s_ready <= emi(13);�   !   #             clk    <= emi(14);�                   emo(10)  <= m_ready;�                   m_last   <= emi(9);5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                            "                    V       ^��     �         #      1   emo(7   downto 0)    <=     s_data(7 downto 0;5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                            "                    V       ^��     �         #      0   emo(7  downto 0)    <=     s_data(7 downto 0;5�_�   o   q           p           ����                                                                                                                                                                                                                                                                                                                                      "          V       ^��    �   !   #   #         clk             <= emi(14);�      !   #         s_ready         <= emi(13);�          #         emo(12)         <= s_last;�         #         emo(11)         <= s_valid;�         #      (   emo(7 downto 0) <= s_data(7 downto 0;�         #         emo(10)         <= m_ready;�         #         m_last          <= emi(9);�         #         m_valid         <= emi(8);�         #      &   m_data          <= emi(7 downto 0);�         #      #           clk     : out STD_LOGIC;�         #      $           s_ready : out STD_LOGIC);�         #      #           s_last  : in  STD_LOGIC;�         #      #           s_valid : in  STD_LOGIC;�         #      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         #      $           m_ready : in  STD_LOGIC);�   
      #      #           m_last  : out STD_LOGIC;�   	      #      #           m_valid : out STD_LOGIC;�      
   #      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   #      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         #      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         #          Port(  �                "   m_data  <=     emi(7 downto 0);�                /   emo(7 downto 0)    <=     s_data(7 downto 0;�                   emo(11) <=     s_valid;�                   m_valid <=     emi(8);�                    emo(12) <=     s_last;�      !             s_ready <=     emi(13);�   !   #             clk     <=     emi(14);�                   emo(10) <=     m_ready;�                   m_last  <=     emi(9);5�_�   p   r           q      "    ����                                                                                                                                                                                                                                                                                                                                      "          V       ^��     �         #      $           s_ready : out STD_LOGIC);5�_�   q   s           r      "    ����                                                                                                                                                                                                                                                                                                                                      "          V       ^��    �         #      #           clk     : out STD_LOGIC;5�_�   r   t           s      "    ����                                                                                                                                                                                                                                                                                                                                      "          V       ^��    �         #      $           m_ready : in  STD_LOGIC);5�_�   s   u           t      '    ����                                                                                                                                                                                                                                                                                                                                      "          V       ^��   	 �         #      (   emo(7 downto 0) <= s_data(7 downto 0;5�_�   t   v           u           ����                                                                                                                                                                                                                                                                                                                                      "          V       ^�~     �         #    �         #    5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                                      #          V       ^�     �         $      $           clk     : out STD_LOGIC);5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                                      #          V       ^��     �         $      %           leds     : out STD_LOGIC);5�_�   w   y           x      "    ����                                                                                                                                                                                                                                                                                                                                      #          V       ^��     �         $      $           leds    : out STD_LOGIC);5�_�   x   z           y      "    ����                                                                                                                                                                                                                                                                                                                                      #          V       ^��     �         $      $           clk     : out STD_LOGIC);5�_�   y   {           z      "    ����                                                                                                                                                                                                                                                                                                                                      #          V       ^��     �         $    5�_�   z   |           {   $       ����                                                                                                                                                                                                                                                                                                                                      $          V       ^��     �   $   '   &         �   $   &   %    5�_�   {   }           |   &   
    ����                                                                                                                                                                                                                                                                                                                                      $          V       ^��     �   %   '   '      
   leds <=5�_�   |   ~           }   &       ����                                                                                                                                                                                                                                                                                                                                      $          V       ^��     �   %   '   '         leds <= 5�_�   }              ~           ����                                                                                                                                                                                                                                                                                                                            &                    V       ^�     �   %   '   '         leds            <=�   #   %   '         clk             <= emi(14);�   !   #   '         s_ready         <= emi(13);�       "   '         emo(12)         <= s_last;�      !   '         emo(11)         <= s_valid;�          '      )   emo(7 downto 0) <= s_data(7 downto 0);�         '         emo(10)         <= m_ready;�         '         m_last          <= emi(9);�         '         m_valid         <= emi(8);�         '      &   m_data          <= emi(7 downto 0);�         '      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         '      #           clk     : out STD_LOGIC;�         '      #           s_ready : out STD_LOGIC;�         '      #           s_last  : in  STD_LOGIC;�         '      #           s_valid : in  STD_LOGIC;�         '      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         '      #           m_ready : in  STD_LOGIC;�   
      '      #           m_last  : out STD_LOGIC;�   	      '      #           m_valid : out STD_LOGIC;�      
   '      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   '      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         '      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         '          Port(  �                &   m_data          <= emi(7 downto 0);�       "             emo(12)         <= s_last;�   %   '             leds <=  �                 )   emo(7 downto 0) <= s_data(7 downto 0);�      !             emo(11)         <= s_valid;�   !   #             s_ready         <= emi(13);�   #   %             clk             <= emi(14);�                   emo(10)         <= m_ready;�                   m_last          <= emi(9);�                   m_valid         <= emi(8);5�_�   ~   �              &       ����                                                                                                                                                                                                                                                                                                                            &                    V       ^�     �   %   '   '         leds            <=5�_�      �           �   &       ����                                                                                                                                                                                                                                                                                                                            &                    V       ^�+     �   %   '   '      )   leds            <= emi( 15 downto 15);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            &                    V       ^�-     �   %   '   '      )   leds            <= emi( 17 downto 15);5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            &                    V       ^�1     �   $   %           5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�>     �   $   &   &      (   leds            <= emi(17 downto 15);5�_�   �   �           �   %   '    ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�@     �   $   &   &      (   leds            <= em9(17 downto 15);5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�J     �   $   &   &      0   leds            <= em9(17 downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�K     �   $   &   &      /   eds            <= em9(17 downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�N     �   $   &   &         em9(17 downto 15) => leds;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�S     �   $   &   &         emi(17 downto 15) => leds;�   #   %   &          clk               <= emi(14);�   !   #   &          s_ready           <= emi(13);�       "   &         emo(12)           <= s_last;�      !   &          emo(11)           <= s_valid;�          &      +   emo(7 downto 0)   <= s_data(7 downto 0);�         &          emo(10)           <= m_ready;�         &         m_last            <= emi(9);�         &         m_valid           <= emi(8);�         &      (   m_data            <= emi(7 downto 0);�         &      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         &      #           clk     : out STD_LOGIC;�         &      #           s_ready : out STD_LOGIC;�         &      #           s_last  : in  STD_LOGIC;�         &      #           s_valid : in  STD_LOGIC;�         &      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         &      #           m_ready : in  STD_LOGIC;�   
      &      #           m_last  : out STD_LOGIC;�   	      &      #           m_valid : out STD_LOGIC;�      
   &      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   &      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         &      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         &          Port(  �                &   m_data          <= emi(7 downto 0);�       "             emo(12)         <= s_last;�   $   &             emi(17 downto 15) => leds;�                 )   emo(7 downto 0) <= s_data(7 downto 0);�      !             emo(11)         <= s_valid;�   !   #             s_ready         <= emi(13);�   #   %             clk             <= emi(14);�                   emo(10)         <= m_ready;�                   m_last          <= emi(9);�                   m_valid         <= emi(8);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�^     �   $   &   &      $   emi(17  downto 15)   =>     leds;�   #   %   &         clk     <=     emi(14);�   !   #   &         s_ready <=     emi(13);�       "   &         emo(12) <=     s_last;�      !   &         emo(11) <=     s_valid;�          &      2   emo(7   downto 0)    <=     s_data(7 downto 0);�         &         emo(10) <=     m_ready;�         &         m_last  <=     emi(9);�         &         m_valid <=     emi(8);�         &      "   m_data  <=     emi(7 downto 0);�         &      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         &      #           clk     : out STD_LOGIC;�         &      #           s_ready : out STD_LOGIC;�         &      #           s_last  : in  STD_LOGIC;�         &      #           s_valid : in  STD_LOGIC;�         &      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         &      #           m_ready : in  STD_LOGIC;�   
      &      #           m_last  : out STD_LOGIC;�   	      &      #           m_valid : out STD_LOGIC;�      
   &      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   &      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         &      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         &          Port(  �       "             emo(12)           <= s_last;�   $   &             emi(17 downto 15) => leds;�                 +   emo(7 downto 0)   <= s_data(7 downto 0);�      !              emo(11)           <= s_valid;�   !   #              s_ready           <= emi(13);�   #   %              clk               <= emi(14);�                    emo(10)           <= m_ready;�                   m_last            <= emi(9);�                   m_valid           <= emi(8);�                (   m_data            <= emi(7 downto 0);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�`     �   $   &   &         emi(17  downto 15) => leds;�   #   %   &      !   clk                <= emi(14);�   !   #   &      !   s_ready            <= emi(13);�       "   &          emo(12)            <= s_last;�      !   &      !   emo(11)            <= s_valid;�          &      ,   emo(7   downto 0)  <= s_data(7 downto 0);�         &      !   emo(10)            <= m_ready;�         &          m_last             <= emi(9);�         &          m_valid            <= emi(8);�         &      )   m_data             <= emi(7 downto 0);�         &      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         &      #           clk     : out STD_LOGIC;�         &      #           s_ready : out STD_LOGIC;�         &      #           s_last  : in  STD_LOGIC;�         &      #           s_valid : in  STD_LOGIC;�         &      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         &      #           m_ready : in  STD_LOGIC;�   
      &      #           m_last  : out STD_LOGIC;�   	      &      #           m_valid : out STD_LOGIC;�      
   &      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   &      8           emo     : out STD_LOGIC_VECTOR (15 downto 0);�         &      8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);�         &          Port(  �                "   m_data  <=     emi(7 downto 0);�       "             emo(12) <=     s_last;�   $   &          $   emi(17  downto 15)   =>     leds;�                 2   emo(7   downto 0)    <=     s_data(7 downto 0);�      !             emo(11) <=     s_valid;�   !   #             s_ready <=     emi(13);�   #   %             clk     <=     emi(14);�                   emo(10) <=     m_ready;�                   m_last  <=     emi(9);�                   m_valid <=     emi(8);5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %                    V       ^�o   
 �   $   &   &         emi(17  downto 15) => leds;5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��     �                8           emi     : in  STD_LOGIC_VECTOR (15 downto 0);5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��    �      	          8           emo     : out STD_LOGIC_VECTOR (15 downto 0);5�_�   �   �           �      6    ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�    �         &      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�H     �   $   &   &         emi(18  downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�I     �   $   &   &         em9(18  downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�J    �   $   &   &         em0(18  downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�g     �   $   &   &         emo(18  downto 15) => leds;5�_�   �   �           �   %   
    ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�i     �   $   &   &      %   leds <=emo(18  downto 15) => leds;5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�l     �   $   &   &      &   leds <= emo(18  downto 15) => leds;5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�o    �   $   &   &      +   leds              <= emo(18  downto 15);�   #   %   &          clk               <= emi(14);�   !   #   &          s_ready           <= emi(13);�       "   &         emo(12)           <= s_last;�      !   &          emo(11)           <= s_valid;�          &      +   emo(7   downto 0) <= s_data(7 downto 0);�         &          emo(10)           <= m_ready;�         &         m_last            <= emi(9);�         &         m_valid           <= emi(8);�         &      (   m_data            <= emi(7 downto 0);�         &      8           leds    : out STD_LOGIC_VECTOR (3 downto 0));�         &      #           clk     : out STD_LOGIC;�         &      #           s_ready : out STD_LOGIC;�         &      #           s_last  : in  STD_LOGIC;�         &      #           s_valid : in  STD_LOGIC;�         &      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         &      #           m_ready : in  STD_LOGIC;�   
      &      #           m_last  : out STD_LOGIC;�   	      &      #           m_valid : out STD_LOGIC;�      
   &      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   &      8           emo     : out STD_LOGIC_VECTOR (31 downto 0);�         &      8           emi     : in  STD_LOGIC_VECTOR (31 downto 0);�         &          Port(  �                )   m_data             <= emi(7 downto 0);�       "              emo(12)            <= s_last;�   $   &             leds <= emo(18  downto 15);�                 ,   emo(7   downto 0)  <= s_data(7 downto 0);�      !          !   emo(11)            <= s_valid;�   !   #          !   s_ready            <= emi(13);�   #   %          !   clk                <= emi(14);�                !   emo(10)            <= m_ready;�                    m_last             <= emi(9);�                    m_valid            <= emi(8);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�z    �   $   &   &      +   leds              <= emo(18  downto 15);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��     �   $   &   &      +   leds              <= emi(18  downto 15);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��     �   $   &   &      +   leds              <= emi(18  downto 15);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��     �   $   &   &      +   leds              <= emi(19  downto 15);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��     �   $   &   &      +   leds              <= emi(18  downto 15);5�_�   �   �           �   %       ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^��    �   $   &   &      +   leds              <= emi(17  downto 15);5�_�   �   �           �          ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�\     �         &      #           clk     : out STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�^     �         &      %           s_clk     : out STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�^     �         &      $           s_clk    : out STD_LOGIC;5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                      %                    V       ^�a     �         &    �         &    5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &                    V       ^�c     �         '      #           s_clk   : out STD_LOGIC;5�_�   �   �           �   %        ����                                                                                                                                                    &                                                                                                                                                                      %          %          V       ^�f     �   $   %              clk               <= emi(14);5�_�   �   �           �          ����                                                                                                                                                    %                                                                                                                                                                      %          %          V       ^�j     �         &    �         &    5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�l     �         '          clk               <= emi(14);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�m     �         '          clk               <= emi(19);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�o     �         '          clk               <= emi(10);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�s     �         '      "   m_clk               <= emi(10);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�s     �         '      !   m_clk              <= emi(10);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                      &          &          V       ^�|     �          '          emo(10)           <= m_ready;5�_�   �   �           �           ����                                                                                                                                                    &                                                                                                                                                                                          V       ^Ҏ     �                    m_clk             <= emi(10);5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                                          V       ^ҏ     �          &    �          &    5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                          V       ^ґ     �         '          emo(11)           <= m_ready;5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                          V       ^Ғ     �         '          emo(19)           <= m_ready;5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                          V       ^ғ     �         '          emo(19)           <= m_ready;5�_�   �   �           �           ����                                                                                                                                                    &                                                                                                                                                                                          V       ^ҕ     �                    m_clk             <= emi(10);5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                                          V       ^Ҙ     �          &    �          &    5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                            V       ^ҟ     �          '          m_clk             <= emi(10);5�_�   �   �           �           ����                                                                                                                                                    &                                                                                                                                                                                          V       ^ҡ     �                    m_clk             <= emi(11);5�_�   �   �           �           ����                                                                                                                                                    %                                                                                                                                                                                          V       ^ҡ     �         &    �         &    5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                            V       ^Ҧ     �         '          m_clk             <= emi(11);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                            V       ^ҧ     �         '          m_clk             <= emi(19);5�_�   �   �           �          ����                                                                                                                                                    &                                                                                                                                                                                            V       ^ҩ     �          '          emo(10)           <= m_ready;5�_�   �   �           �   "       ����                                                                                                                                                    &                                                                                                                                                                                            V       ^Ү     �   !   #   '          emo(11)           <= s_valid;5�_�   �   �           �   #       ����                                                                                                                                                    &                                                                                                                                                                                            V       ^Ү     �   "   $   '         emo(12)           <= s_last;5�_�   �   �           �   $       ����                                                                                                                                                    &                                                                                                                                                                                            V       ^Ҳ     �   #   %   '    �   $   %   '    5�_�   �   �           �   $       ����                                                                                                                                                    '                                                                                                                                                                                            V       ^ҵ     �   #   %   (          m_clk             <= emi(10);5�_�   �   �           �   $       ����                                                                                                                                                    '                                                                                                                                                                                            V       ^ҷ     �   #   %   (          s_clk             <= emi(10);5�_�   �   �           �   $       ����                                                                                                                                                    '                                                                                                                                                                                            V       ^Ҹ     �   #   %   (          s_clk             <= emi(13);5�_�   �   �           �   %       ����                                                                                                                                                    '                                                                                                                                                                                            V       ^Һ     �   $   &   (          s_ready           <= emi(13);5�_�   �   �           �   '   2    ����                                                                                                                                                    '                                                                                                                                                                                            V       ^��     �   &   (   (      5   leds              <= emi(13) & emi(17  downto 15);5�_�   �   �           �   '   '    ����                                                                                                                                                    '                                                                                                                                                                                            V       ^��     �   &   (   (      5   leds              <= emi(13) & emi(17  downto 16);5�_�   �   �           �   '       ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^��     �   &   (   (      5   leds              <= emi(13) & emi(18  downto 16);5�_�   �   �           �   '       ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^��    �   &   (   (      +   leds              <= emi(18  downto 16);5�_�   �   �           �   '       ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^��     �   &   (   (      +   leds              <= emi(19  downto 16);5�_�   �   �           �   '   -    ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^��    �   &   (   (      ;   leds              <= s_clk & m_clk & emi(19  downto 16);5�_�   �   �           �   '   -    ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^�W     �   '   )   )         �   '   )   (    5�_�   �   �           �           ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^�p     �         )    �         )    5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�q     �         *      #           s_clk   : out STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�r     �         *      !           rst   : out STD_LOGIC;5�_�   �   �           �      6    ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�u     �         *      8           leds    : out STD_LOGIC_VECTOR (3 downto 0));5�_�   �   �           �      "    ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�v    �         *      #           rst     : out STD_LOGIC;5�_�   �   �           �   )       ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^��    �   (   *   *         rst               <= emi(20)5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�8     �         *      $           rst     : out STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�9     �         *      %           rsto     : out STD_LOGIC);5�_�   �   �           �   )       ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�<     �   (   *   *          rst               <= emi(20);5�_�   �   �           �   )       ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�=    �   (   *   *      !   rsto               <= emi(20);5�_�   �   �           �   )       ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�     �   (   )              rsto              <= emi(20);5�_�   �   �           �      
    ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�     �                $           rsto    : out STD_LOGIC);5�_�   �   �           �      6    ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^�    �         (      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);5�_�   �   �           �           ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^�%     �         (       5�_�   �   �           �          ����                                                                                                                                                    '                                                                                                                                                                      '          '   !       v   !    ^�=     �         (    �         (    5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�?     �         )      signal s_clk_sig: STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�?     �         )      signal m_clk_sig: STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�@     �         )      signal ,_clk_sig: STD_LOGIC;5�_�   �   �           �   &       ����                                                                                                                                                    (                                                                                                                                                                      (          (   !       v   !    ^�G     �   &   (   )    �   &   '   )    5�_�   �   �           �   '        ����                                                                                                                                                    )                                                                                                                                                                      '           '          v       ^�I     �   &   (   *      signal s_clk_sig: STD_LOGIC;5�_�   �   �           �   '        ����                                                                                                                                                    )                                                                                                                                                                      '           '          v       ^�K     �   &   (   *      s_clk_sig: STD_LOGIC;5�_�   �   �           �   '       ����                                                                                                                                                    )                                                                                                                                                                      '           '          v       ^�L     �   &   (   *         s_clk_sig: STD_LOGIC;5�_�   �   �           �   '       ����                                                                                                                                                    )                                                                                                                                                                      '          '          v       ^�R     �   &   (   *         s_clk_sig <= : STD_LOGIC;5�_�   �   �           �   '       ����                                                                                                                                                    )                                                                                                                                                                      '          '          v       ^�W     �   &   (   *         s_clk_sig <= clk;5�_�   �   �           �   )       ����                                                                                                                                                    )                                                                                                                                                                      '          '          v       ^�\     �   (   *   *      ;   leds              <= s_clk & m_clk & emi(17  downto 16);5�_�   �   �           �   '       ����                                                                                                                                                    )                                                                                                                                                                      '          '          v       ^�_     �   &   (   +         �   &   (   *    5�_�   �   �           �   (       ����                                                                                                                                                    *                                                                                                                                                                      (          (          v       ^�a     �   '   )   +    �   (   )   +    5�_�   �   �           �   )       ����                                                                                                                                                    +                                                                                                                                                                      )          )          v       ^�c     �   (   *   ,         s_clk_sig <= s_clk;5�_�   �   �           �   )       ����                                                                                                                                                    +                                                                                                                                                                      )          )          v       ^�d     �   (   *   ,         m_clk_sig <= s_clk;5�_�   �   �           �   '       ����                                                                                                                                                    +                                                                                                                                                                      )          )          v       ^�e     �   &   '             P5�_�   �   �           �   *   )    ����                                                                                                                                                    *                                                                                                                                                                      (          (          v       ^�g     �   )   +   +      ?   leds              <= s_clk_sig & m_clk & emi(17  downto 16);5�_�   �   �           �           ����                                                                                                                                                    *                                                                                                                                                                                          V   ,    ^�n    �                signal m_clk_sig: STD_LOGIC;�                signal s_clk_sig: STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    *                                                                                                                                                                                          V   ,    ^�     �         +    �         +    5�_�   �   �           �      "    ����                                                                                                                                                    +                                                                                                                                                                                          V   ,    ^�     �         ,      #           s_clk   : out STD_LOGIC;5�_�   �   �           �      6    ����                                                                                                                                                    +                                                                                                                                                                                          V   ,    ^�     �         ,      8           leds    : out STD_LOGIC_VECTOR (3 downto 0));5�_�   �   �           �          ����                                                                                                                                                    +                                                                                                                                                                                          V   ,    ^�     �         ,      $           s_clk   : out STD_LOGIC);5�_�   �   �   �       �   )       ����                                                                                                                                                    +                                                                                                                                                                                          V   ,    ^�     �   (   *   ,    �   )   *   ,    5�_�   �   �           �   *       ����                                                                                                                                                    ,                                                                                                                                                                      *          *          v       ^�     �   )   +   -         m_clk_sig <= m_clk;5�_�   �   �           �   *   
    ����                                                                                                                                                    ,                                                                                                                                                                      *          *          v       ^�     �   )   +   -         rst <= m_clk;5�_�   �   �           �   *   
    ����                                                                                                                                                    ,                                                                                                                                                                      '          '          v       ^�     �   )   +   -         rst <= ;�   *   +   -    5�_�   �   �           �   *       ����                                                                                                                                                    ,                                                                                                                                                                      '          '          v       ^�    �   )   *             rst <= emi(15);5�_�   �   �           �          ����                                                                                                                                                    +                                                                                                                                                                                                 ^��    �         ,         signal m_clk_sig: STD_LOGIC;�         ,         signal s_clk_sig: STD_LOGIC;5�_�   �   �           �   )       ����                                                                                                                                                    +                                                                                                                                                                                                 ^��     �   (   *   ,    �   )   *   ,    5�_�   �   �           �   *       ����                                                                                                                                                    ,                                                                                                                                                                                                 ^��     �   )   +   -         m_clk_sig <= m_clk;5�_�   �   �           �   *   
    ����                                                                                                                                                    ,                                                                                                                                                                                                 ^��    �   )   +   -         tst <= m_clk;5�_�   �   �           �   *       ����                                                                                                                                                    ,                                                                                                                                                                                                 ^��    �   )   +   -         tst <= emi(20);5�_�   �   �           �          ����                                                                                                                                                    ,                                                                                                                                                                                                 ^�    �         -      %   signal s_clk_sig: inout STD_LOGIC;   %   signal m_clk_sig: inout STD_LOGIC;5�_�   �   �           �   ,       ����                                                                                                                                                    ,                                                                                                                                                                                                 ^�>     �   +   -   -    �   ,   -   -    5�_�   �   �           �   -       ����                                                                                                                                                    -                                                                                                                                                                      -          -   /       v   /    ^�A     �   ,   .   .      C   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�   �   �           �   -       ����                                                                                                                                                    -                                                                                                                                                                      -          -   /       v   /    ^�C     �   ,   .   .      +   leds              <= emi(17  downto 16);5�_�   �   �           �   ,        ����                                                                                                                                                    -                                                                                                                                                                      -          -   /       v   /    ^�E     �   +   -   .      C   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�   �   �           �   ,        ����                                                                                                                                                    -                                                                                                                                                                      ,           ,                 ^�J    �   +   -   .      E//   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�   �   �           �          ����                                                                                                                                                    -                                                                                                                                                                      ,           ,                 ^�     �         .      #           s_clk   : out STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                    -                                                                                                                                                                      ,           ,                 ^�     �         .      #           m_clk   : out STD_LOGIC;5�_�   �   �           �           ����                                                                                                                                                    -                                                                                                                                                                                          V       ^��     �                   signal s_clk_sig: STD_LOGIC;      signal m_clk_sig: STD_LOGIC;5�_�   �   �           �   '        ����                                                                                                                                                    +                                                                                                                                                                      &           '           V        ^��     �   %   '   +         s_clk_sig <= s_clk;�   &   '             m_clk_sig <= m_clk;5�_�   �   �           �   &       ����                                                                                                                                                    *                                                                                                                                                                      &           '           V        ^��     �   %   &             jjj5�_�   �              �   (        ����                                                                                                                                                    )                                                                                                                                                                      &           &           V        ^��     �   '   )   *      E--   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�   �                (        ����                                                                                                                                                    )                                                                                                                                                                      &           &           V        ^��     �   '   )   *      D-   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�                  (       ����                                                                                                                                                    )                                                                                                                                                                      (          (           v        ^��     �   '   )   *      C   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�                 (   %    ����                                                                                                                                                    )                                                                                                                                                                      (   %       (   (       v   (    ^��     �   '   )   *      ?   leds              <= s_clk & m_clk_sig & emi(17  downto 16);5�_�                 )       ����                                                                                                                                                    )                                                                                                                                                                      (   %       (   (       v   (    ^��    �   (   )          +   leds              <= emi(19  downto 16);5�_�                        ����                                                                                                                                                                                                                                                                                                                           (   %       (   (       v   (    ^�A     �         )      %           s_clk   : inout STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                           (   %       (   (       v   (    ^�A     �         )      $           s_clk   : nout STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                           (   %       (   (       v   (    ^�B     �         )      %           m_clk   : inout STD_LOGIC;5�_�    	                    ����                                                                                                                                                                                                                                                                                                                           (   %       (   (       v   (    ^�C     �         )      $           m_clk   : nout STD_LOGIC;5�_�    
        	   &       ����                                                                                                                                                                                                                                                                                                                           (   %       (   (       v   (    ^�l     �   &   *   *         �   &   (   )    5�_�  	            
   '   
    ����                                                                                                                                                                                                                                                                                                                           +   %       +   (       v   (    ^�x     �   &   (   ,         process 5�_�  
               (       ����                                                                                                                                                                                                                                                                                                                           +   %       +   (       v   (    ^�}     �   (   *   ,    5�_�                        ����                                                                                                                                                                                                                                                                                                                           ,   %       ,   (       v   (    ^�     �         .         �         -    5�_�                        ����                                                                                                                                                                                                                                                                                                                           -   %       -   (       v   (    ^�     �         .    �         .    5�_�                    
    ����                                                                                                                                                                                                                                                                                                                           .   %       .   (       v   (    ^�     �         /         signal s_clk: STD_LOGIC;5�_�                 *       ����                                                                                                                                                                                                                                                                                                                           .   %       .   (       v   (    ^�     �   *   ,   0            �   *   ,   /    5�_�                 +       ����                                                                                                                                                                                                                                                                                                                           /   %       /   (       v   (    ^�     �   +   -   1            �   +   -   0    5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                           0   %       0   (       v   (    ^�     �   +   -   1         end process5�_�                        ����                                                                                                                                                                                                                                                                                                                                                      ^�     �         1         signal m_clk: STD_LOGIC;�         1         signal s_clk: STD_LOGIC;5�_�                 )        ����                                                                                                                                                                                                                                                                                                                           )          ,          V       ^�     �   (   -   1    �   )   *   1    5�_�                 -       ����                                                                                                                                                                                                                                                                                                                           -          0          V       ^�     �   ,   .   5         process (s_clk) 5�_�                 /       ����                                                                                                                                                                                                                                                                                                                           -          0          V       ^�     �   .   0   5            s_clk_sig <= s_clk;5�_�                 /       ����                                                                /                                                                                                                                             /                                                                                                          -          0          V       ^�     �   .   0   5            n_clk_sig <= s_clk;5�_�                 /       ����                                                                /                                                                                                                                             /                                                                                                          -          0          V       ^�     �   .   0   5            _clk_sig <= s_clk;5�_�                 /       ����                                                                /                                                                                                                                             /                                                                                                          -          0          V       ^��     �   .   0   5            m_clk_sig <= s_clk;5�_�                 4       ����                                                                /                                                                                                                                             /                                                                                                          -          0          V       ^��     �   3   5   5      ;   leds              <= s_clk & m_clk & emi(17  downto 16);5�_�                 4   )    ����                                                                /                                                                                                                                             /                                                                                                          -          0          V       ^��    �   3   5   5      ?   leds              <= s_clk_sig & m_clk & emi(17  downto 16);5�_�                 1        ����                                                                /                                                                                                                                             /                                                                                                          1           2          V   ,    ^��     �   0   1                    5�_�                         ����                                                                /                                                                                                                                             /                                                                                                          1           1          V   ,    ^�+     �      !   3    �       !   3    5�_�                 !       ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�-     �       "   4          m_clk             <= emi(10);5�_�                 !       ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�0     �       !          #   m_clk_in             <= emi(10);5�_�                         ����                                                                /                                                                                                                                             /                                                                                                          1           1          V   ,    ^�4     �         3    �         3    5�_�    !                     ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�6     �         4      #           m_clk   : out STD_LOGIC;5�_�     "          !          ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�7     �         4      &           m_clk_in   : out STD_LOGIC;5�_�  !  #          "          ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�7     �         4      %           m_clk_in  : out STD_LOGIC;5�_�  "  $          #          ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�8     �         4      $           m_clk_in : out STD_LOGIC;5�_�  #  &          $          ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�:     �         4    �         4    5�_�  $  '  %      &          ����                                                                1                                                                                                                                             1                                                                                                          3           3          V   ,    ^�=     �         5      #           s_clk   : out STD_LOGIC;5�_�  &  (          '          ����                                                                1                                                                                                                                             1                                                                                                          3           3          V   ,    ^�@     �         5      &           s_clk_in   : out STD_LOGIC;5�_�  '  )          (          ����                                                                1                                                                                                                                             1                                                                                                          3           3          V   ,    ^�A     �         5      %           s_clk_in  : out STD_LOGIC;5�_�  (  *          )          ����                                                                1                                                                                                                                             1                                                                                                          3           3          V   ,    ^�A     �         5      $           s_clk_in : out STD_LOGIC;5�_�  )  +          *           ����                                                                1                                                                                                                                             1                                                                                                                              V       ^�F     �                   signal s_clk_sig: STD_LOGIC;      signal m_clk_sig: STD_LOGIC;5�_�  *  ,          +   )        ����                                                                /                                                                                                                                             /                                                                                                          )           0           V        ^�I     �   (   )             process (s_clk)       begin         s_clk_sig <= s_clk;      end process;      process (m_clk)       begin         m_clk_sig <= m_clk;      end process;5�_�  +  -          ,   *       ����                                                                                                                                                                                                                                                                                                                         )           )           V        ^�M     �   )   +   +      C   leds              <= s_clk_sig & m_clk_sig & emi(17  downto 16);5�_�  ,  .          -   *   (    ����                                                                                                                                                                                                                                                                                                                         )           )           V        ^�O     �   )   +   +      B   leds              <= s_clk_in & m_clk_sig & emi(17  downto 16);5�_�  -  /          .   *   (    ����                                                                                                                                                                                                                                                                                                                         )           )           V        ^�Q   ! �   )   +   +      @   leds              <= s_clk_in & m_clkin & emi(17  downto 16);5�_�  .  0          /   #        ����                                                                                                                                                                                                                                                                                                                         (          #   "       V   "    ^�   " �   )   +   +      A   leds              <= s_clk_in & m_clk_in & emi(17  downto 16);�   '   )   +          rst               <= emi(20);�   &   (   +          s_ready           <= emi(15);�   %   '   +          s_clk             <= emi(14);�   $   &   +         emo(13)           <= s_last;�   #   %   +          emo(12)           <= s_valid;�   "   $   +      +   emo(7   downto 0) <= s_data(7 downto 0);�       "   +          emo(11)           <= m_ready;�      !   +          m_clk             <= emi(10);�          +         m_last            <= emi(9);�         +         m_valid           <= emi(8);�         +      (   m_data            <= emi(7 downto 0);�         +      "           rst   : out STD_LOGIC);�         +      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         +      #           s_clk_in : in STD_LOGIC;�         +      #           s_clk   : out STD_LOGIC;�         +      #           s_ready : out STD_LOGIC;�         +      #           s_last  : in  STD_LOGIC;�         +      #           s_valid : in  STD_LOGIC;�         +      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         +      #           m_clk_in : in STD_LOGIC;�         +      #           m_clk   : out STD_LOGIC;�         +      #           m_ready : in  STD_LOGIC;�   
      +      #           m_last  : out STD_LOGIC;�   	      +      #           m_valid : out STD_LOGIC;�      
   +      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   +      8           emo     : out STD_LOGIC_VECTOR (31 downto 0);�         +      8           emi     : in  STD_LOGIC_VECTOR (31 downto 0);�         +          Port(  �   "   $          +   emo(7   downto 0) <= s_data(7 downto 0);�   '   )             rst <= emi(20);�   &   (              s_ready           <= emi(15);�   %   '              s_clk             <= emi(14);�   $   &             emo(13)           <= s_last;�   #   %              emo(12)           <= s_valid;5�_�  /  1          0           ����                                                                                                                                                                                                                                                                                                                         (          #   "       V   "    ^�     �          ,         �         +    5�_�  0  2          1           ����                                                                                                                                                                                                                                                                                                                         +          &   "       V   "    ^�     �         .       5�_�  1  3          2          ����                                                                                                                                                                                                                                                                                                                         +          &   "       V   "    ^��     �      !   .         one_shot:process(5�_�  2  4          3          ����                                                                                                                                                                                                                                                                                                                         -          (   "       V   "    ^��     �      "   1            �      !   0    5�_�  3  5          4   !        ����                                                                                                                                                                                                                                                                                                                         /          *   "       V   "    ^��     �       !          begin5�_�  4  6          5           ����                                                                                                                                                                                                                                                                                                                         .          )   "       V   "    ^��     �       "   2      	         �       "   1    5�_�  5  7          6            ����                                                                                                                                                                                                                                                                                                                         /          *   "       V   "    ^��     �       "   3      	         �       "   2    5�_�  6  8          7           ����                                                                                                                                                                                                                                                                                                                         0          +   "       V   "    ^��     �       "   3    5�_�  7  9          8   "   	    ����                                                                                                                                                                                                                                                                                                                         1          ,   "       V   "    ^��     �   !   #   4               end if;5�_�  8  :          9   !        ����                                                                                                                                                                                                                                                                                                                         1          ,   "       V   "    ^��     �       "   4       5�_�  9  ;          :          ����                                                                                                                                                                                                                                                                                                                         1          ,   "       V   "    ^��     �         4         one_shot:process(emi(8)) is:5�_�  :  <          ;           ����                                                                                                                                                                                                                                                                                                                         1          ,   "       V   "    ^��     �      !   4    �       !   4    5�_�  ;  =          <           ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^��     �      !   5      !      if rising_edge(emi(8)) then5�_�  <  >          =           ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^��     �      !   5      #      if rising_edge(m_clk(8)) then5�_�  =  ?          >           ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^��     �      !   5      "      if rising_edge(m_clk8)) then5�_�  >  @          ?           ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^��     �      !   5      !      if rising_edge(m_clk)) then5�_�  ?  A          @   !       ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^��     �       "   5      !      if rising_edge(emi(8)) then5�_�  @  B          A          ����                                                                                                                                                                                                                                                                                                                         2          -   "       V   "    ^�<     �          6            �          5    5�_�  A  C          B      '    ����                                                                                                                                                                                                                                                                                                                         3          .   "       V   "    ^�S     �          6      )      signal last_m_valid: STD_LOGIC :=0;5�_�  B  D          C      )    ����                                                                                                                                                                                                                                                                                                                         3          .   "       V   "    ^�W     �          6      *      signal last_m_valid: STD_LOGIC :='0;5�_�  C  E          D          ����                                                                                                                                                                                                                                                                                                                                             v       ^�^     �          6      +      signal last_m_valid: STD_LOGIC :='0';5�_�  D  F          E          ����                                                                                                                                                                                                                                                                                                                                             v       ^�n     �         6      %   one_shot:process(m_clk,emi(8)) is:5�_�  E  G          F   "       ����                                                                                                                                                                                                                                                                                                                                             v       ^�u     �   !   $   6      $         if rising_edge(emi(8)) then5�_�  F  H          G   "       ����                                                                                                                                                                                                                                                                                                                                             v       ^��     �   !   #   7      2         if last_m_valid = '0' and emi(8)='1' then5�_�  G  I          H   "   .    ����                                                                                                                                                                                                                                                                                                                                             v       ^��     �   !   #   7      3         if (last_m_valid = '0' and emi(8)='1' then5�_�  H  J          I   #       ����                                                                                                                                                                                                                                                                                                                                             v       ^��     �   "   $   7      $            rising_edge(emi(8)) then5�_�  I  K          J   #       ����                                                                                                                                                                                                                                                                                                                         #          #   2       v   2    ^��     �   "   $   7      3            m_valid <= '1'lrising_edge(emi(8)) then5�_�  J  M          K   "       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   !   #   7      4         if (last_m_valid = '0' and emi(8)='1') then5�_�  K  N  L      M   $       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   #   %   7      	         �   $   %   7    5�_�  M  O          N   $       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   #   %                  last_m_valid 5�_�  N  P          O   $       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   #   %   7                  last_m_valid 5�_�  O  Q          P   $       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   $   &   8                  �   $   &   7    5�_�  P  R          Q   %   	    ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   $   &   8               end if;5�_�  Q  S          R   "       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   !   $   8      4         if (last_m_valid = '0' and emi(8)='1') then5�_�  R  T          S   #   	    ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�      �   "   $   9      !         if( and emi(8)='1') then5�_�  S  U          T   "        ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�     �   !   #   9                if (last_m_valid = '0')5�_�  T  V          U   &   	    ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�     �   %   '   9                  else end if;5�_�  U  W          V   &   	    ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�     �   %   '   9                 else end if;5�_�  V  X          W   &   	    ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�     �   %   '   9                else end if;5�_�  W  Y          X   &       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^�	     �   %   (   9               else end if;5�_�  X  Z          Y   #       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�     �   "   $   :      $            if( and emi(8)='1') then5�_�  Y  [          Z   #       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�!     �   "   $   :      $            if( lnd emi(8)='1') then5�_�  Z  \          [   $       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�&     �   #   %                      m_valid <= '1';5�_�  [  ]          \   %       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�+     �   $   &          !            last_m_valid := '1'; 5�_�  \  ^          ]   &       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�1     �   &   (   :    5�_�  ]  _          ^   '        ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�2     �   '   )   ;    �   '   (   ;    5�_�  ^  `          _   '        ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�3     �   &   '           5�_�  _  a          `   '       ����                                                                                                                                                                                                                                                                                                                         #          #          v       ^�4     �   &   (   ;                     m_valid <= '1';5�_�  `  b          a   $        ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^�W     �   9   ;   ;      A   leds              <= s_clk_in & m_clk_in & emi(17  downto 16);�   7   9   ;          rst               <= emi(20);�   6   8   ;          s_ready           <= emi(15);�   5   7   ;          s_clk             <= emi(14);�   4   6   ;         emo(13)           <= s_last;�   3   5   ;          emo(12)           <= s_valid;�   2   4   ;      +   emo(7   downto 0) <= s_data(7 downto 0);�   0   2   ;          emo(11)           <= m_ready;�   /   1   ;          m_clk             <= emi(10);�   .   0   ;         m_last            <= emi(9);�   -   /   ;         m_valid           <= emi(8);�   ,   .   ;      (   m_data            <= emi(7 downto 0);�   *   ,   ;         end process one_shot;�   )   +   ;      	         �   (   *   ;            end if;�   '   )   ;               end if;�   &   (   ;                     m_valid <= '0';�   %   '   ;               else �   $   &   ;      #               last_m_valid := '1';�   #   %   ;      #               m_valid      <= '1';�   "   $   ;                  if(emi(8)='1') then�   !   #   ;      %         if (last_m_valid = '0') then�       "   ;             if rising_edge(m_clk) then�      !   ;         begin�          ;      -      variable last_m_valid: STD_LOGIC :='0';�         ;         one_shot:process(m_clk) is:�         ;      "           rst   : out STD_LOGIC);�         ;      7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�         ;      #           s_clk_in : in STD_LOGIC;�         ;      #           s_clk   : out STD_LOGIC;�         ;      #           s_ready : out STD_LOGIC;�         ;      #           s_last  : in  STD_LOGIC;�         ;      #           s_valid : in  STD_LOGIC;�         ;      8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);�         ;      #           m_clk_in : in STD_LOGIC;�         ;      #           m_clk   : out STD_LOGIC;�         ;      #           m_ready : in  STD_LOGIC;�   
      ;      #           m_last  : out STD_LOGIC;�   	      ;      #           m_valid : out STD_LOGIC;�      
   ;      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);�      	   ;      8           emo     : out STD_LOGIC_VECTOR (31 downto 0);�         ;      8           emi     : in  STD_LOGIC_VECTOR (31 downto 0);�         ;          Port(  �   #   %                         m_valid <= '1';�   $   &          $               last_m_valid := '1'; 5�_�  a  c          b   (       ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^�^     �   '   )   ;    �   (   )   ;    5�_�  b  d          c   %        ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^�j     �   %   '   =                     �   %   '   <    5�_�  c  e          d   )       ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^��     �   (   +   =      #               last_m_valid := '1';5�_�  d  f          e   )       ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^��     �   (   *   >                     if(emi(8)='0')5�_�  e  g          f   *        ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^��     �   )   +   >      #               last_m_valid := '1';5�_�  f  h          g   *        ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^��     �   *   ,   ?                     �   *   ,   >    5�_�  g  i          h   *       ����                                                                                                                                                                                                                                                                                                                         $          %          V       ^��     �   )   +          #               last_m_valid := '0';5�_�  h  j          i   (        ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �   )   +          &                  last_m_valid := '0';�   (   *          "               if(emi(8)='0') then�   '   )                         m_valid <= '0';5�_�  i  k          j   .       ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �   -   .          	         5�_�  j  l          k          ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��   # �          >      -      variable last_m_valid: STD_LOGIC :='0';5�_�  k  m          l   %       ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �   $   &   >      #               last_m_valid := '1';5�_�  l  n          m   %       ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �   $   &   >      #               last_m_valid >= '1';5�_�  m  o          n   *       ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �   )   +   >      #               last_m_valid := '0';5�_�  n  p          o   1       ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^�Q   $ �   0   2   >         m_valid           <= emi(8);5�_�  o  q          p          ����                                                                                                                                                                                                                                                                                                                         (          +          V       ^��     �         >         one_shot:process(m_clk) is:5�_�  p  r          q          ����                                                                                                                                                                                                                                                                                                                                             v       ^��     �         >      $   one_shot:process(emi(10m_clk) is:5�_�  q  s          r          ����                                                                                                                                                                                                                                                                                                                                             v       ^��   % �         >         one_shot:process(emi(10) is:5�_�  r  t          s          ����                                                                                                                                                                                                                                                                                                                                             v       ^��   & �         >          one_shot:process(emi(10)) is:5�_�  s  u          t           ����                                                                                                                                                                                                                                                                                                                                               V        ^��     �                +      signal last_m_valid: STD_LOGIC :='0';5�_�  t  v          u          ����                                                                                                                                                                                                                                                                                                                                               V        ^�   ' �         =    �         =    5�_�  u  w          v   !       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�   ( �       "   >             if rising_edge(m_clk) then5�_�  v  x          w          ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�W     �          >         one_shot:process(emi(10)) is5�_�  w  y          x           ����                                                                                                                                                                                                                                                                                                                                   .          V       ^�`     �      /   >    �          >    5�_�  x  z          y   .       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�c     �   -   /   N         end process one_shot;5�_�  y  {          z   /       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�g     �   .   0   N      !   m_one_shot:process(emi(10)) is5�_�  z  |          {   >       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�j     �   =   ?   N         end process one_shot;5�_�  {  }          |   >       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�l     �   =   ?   N         end process s)one_shot;5�_�  |  ~          }   >       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�m     �   =   ?   N         end process s)one_shot;5�_�  }            ~   .       ����                                                                                                                                                                                                                                                                                                                         /          >          V       ^�r     �   .   0   N    5�_�  ~  �                     ����                                                                                                                                                                                                                                                                                                                         0          ?          V       ^��     �         O    �         O    5�_�    �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P      #           s_clk_in : in STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P      "           _clk_in : in STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P      !           clk_in : in STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P                  clkin : in STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P                 clkn : in STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         1          @          V       ^��     �         P                 clk : in STD_LOGIC;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �      !   P      !   m_one_shot:process(emi(10)) is5�_�  �  �          �   "       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   !   #   P      "      if rising_edge(emi(10)) then5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   2   4   P      "      if rising_edge(emi(10)) then5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   0   2   P      !   s_one_shot:process(emi(10)) is5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   3   5   P      %         if (last_m_valid = '0') then5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   3   5   P      %         if (last_s_valid = '0') then5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �   K   M   P          s_ready           <= emi(15);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                               v       ^��     �         P    �         P    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^��     �         Q      +      signal last_m_valid: STD_LOGIC :='0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^��     �         Q      +      signal last_s_valid: STD_LOGIC :='0';5�_�  �  �          �   6       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   5   7   Q                  if(emi(8)='1') then5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   6   8   Q      #               m_valid      <= '1';5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   6   8   Q      #               s_valid      <= '1';5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   7   9   Q      #               last_m_valid <= '1';5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   7   9   Q      #               last_s_valid <= '1';5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   :   <   Q                  m_valid <= '0';5�_�  �  �          �   ;       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   :   <   Q                  s_valid <= '0';5�_�  �  �          �   <       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   ;   =   Q                  if(emi(8)='0') then5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�     �   <   >   Q      #               last_m_valid <= '0';5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                         !          !          v       ^�   ) �   <   >   Q      #               last_s_valid <= '0';5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                               V        ^�     �                #           m_clk   : out STD_LOGIC;   #           m_clk_in : in STD_LOGIC;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                               V        ^�     �                #           s_clk   : out STD_LOGIC;   #           s_clk_in : in STD_LOGIC;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                               V        ^�0     �         M    �         M    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                               V        ^�A     �         N         m_one_shot:process(clk) is5�_�  �  �  �      �      
    ����                                                                                                                                                                                                                                                                                                                                               V        ^�J     �         O            �         N    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                               V        ^�_     �         O    �         O    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                               V        ^�`     �         P            if rst='0' then5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                                               V        ^��     �   "   $   P    �   #   $   P    5�_�  �  �          �   #       ����                                                                                                                                                                                                                                                                                                                                               V        ^��     �   "   %   Q               if rst='0' then5�_�  �  �  �      �   $       ����                                                                                                                                                                                                                                                                                                                                             V       ^��     �   #   %   R    �   $   %   R    5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                                             V       ^��     �   #   %   S      +      signal last_m_valid: STD_LOGIC :='0';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                         $          $          v       ^��     �   #   %   S      1            signal last_m_valid: STD_LOGIC :='0';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                         $          $          v       ^��     �   #   %   S      *            last_m_valid: STD_LOGIC :='0';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                         $          $   )       v   )    ^��     �   #   %   S      -            last_m_valid <=: STD_LOGIC :='0';5�_�  �  �          �   %       ����                                                                                                                                                                                                                                                                                                                         $          $   )       v   )    ^��     �   $   &   S                  5�_�  �  �          �   &        ����                                                                                                                                                                                                                                                                                                                         &   	       0   	       V   	    ^��     �   /   1                   end if;�   .   0                      end if;�   -   /          #               last_m_valid <= '0';�   ,   .                      if(emi(8)='0') then�   +   -                      m_valid <= '0';�   *   ,                   else �   )   +                      end if;�   (   *          #               last_m_valid <= '1';�   '   )          #               m_valid      <= '1';�   &   (                      if(emi(8)='1') then�   %   '          %         if (last_m_valid = '0') then5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                         &   	       0   	       V   	    ^��     �   /   1   S    �   0   1   S    5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                         &   	       1   	       V   	    ^��     �   0   2                      end if;5�_�  �  �          �   8        ����                                                                                                                                                                                                                                                                                                                         #   	       %   	       V   	    ^��     �   7   ;   T    �   8   9   T    5�_�  �  �  �      �   9       ����                                                                                                                                                                                                                                                                                                                         #   	       %   	       V   	    ^��     �   8   :   W                  last_m_valid <=0';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                         #   	       %   	       V   	    ^��     �   8   :   W                  last_s_valid <=0';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                         #   	       %   	       V   	    ^��     �   8   :   W                  last_s_readyy <=0';5�_�  �  �          �   ;        ����                                                                                                                                                                                                                                                                                                                         ;          E          V       ^��     �   D   F                   end if;�   C   E                      end if;�   B   D          #               last_s_ready <= '0';�   A   C                       if(emi(15)='0') then�   @   B                      s_ready <= '0';�   ?   A                   else �   >   @                      end if;�   =   ?          #               last_s_ready <= '1';�   <   >          #               s_ready      <= '1';�   ;   =                       if(emi(15)='1') then�   :   <          %         if (last_s_ready = '0') then5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                         ;          E          V       ^��     �   D   F   W    �   E   F   W    5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �   E   G                      end if;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �         X      "           rst   : out STD_LOGIC);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �         X      #           rst    : out STD_LOGIC);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �         X      "           rst    : in STD_LOGIC);5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �   L   M              m_clk             <= emi(10);5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                         ;          F          V       ^��     �   Q   R              s_clk             <= emi(14);5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^��     �   T   V   V      A   leds              <= s_clk_in & m_clk_in & emi(17  downto 16);5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^��     �   L   N   V          emo(11)           <= m_ready;5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^��     �   L   N   V          emo(19)           <= m_ready;5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^��     �   O   Q   V          emo(12)           <= s_valid;5�_�  �  �          �   Q       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^�      �   P   R   V         emo(13)           <= s_last;5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^�     �   Q   S   V      "   --s_ready           <= emi(15);5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^�     �   Q   S   V      "   --s_ready           <= emi(14);5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                         U          U   -       v   -    ^�     �   R   S              rst               <= emi(20);5�_�  �  �          �   T   (    ����                                                                                                                                                                                                                                                                                                                         T          T   -       v   -    ^�     �   S   U   U      +   leds              <= emi(17  downto 16);5�_�  �  �          �   <        ����                                                                                                                                                                                                                                                                                                                         :          B          V       ^�(   * �   A   C          #               if(emi(15)='0') then�   ;   =          #               if(emi(15)='1') then5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                         :          B          V       ^�O   + �   #   %   U                  last_m_valid <=0';5�_�  �  �  �      �   9       ����                                                                                                                                                                                                                                                                                                                         :          B          V       ^�Y   , �   8   :   U                  last_s_ready <=0';5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                              V       ^�o     �                   rst_proc:process(clk) is         if rising_edge(clk) then            if rst='0' then    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                              V       ^�p   - �         Q    5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                              V       ^��   . �                 5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         Q      #           m_valid : out STD_LOGIC;   #           m_last  : out STD_LOGIC;   #           m_ready : in  STD_LOGIC;       8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);   #           s_valid : in  STD_LOGIC;   #           s_last  : in  STD_LOGIC;   #           s_ready : out STD_LOGIC;�      	   Q      8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       ^�   / �         Q   	   <           axi)m_data  : out STD_LOGIC_VECTOR (7  downto 0);   '           axi)m_valid : out STD_LOGIC;   '           axi)m_last  : out STD_LOGIC;   '           axi)m_ready : in  STD_LOGIC;       <           axi)s_data  : in  STD_LOGIC_VECTOR (7  downto 0);   '           axi)s_valid : in  STD_LOGIC;   '           axi)s_last  : in  STD_LOGIC;   '           axi)s_ready : out STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       ^�   0 �         Q      '           axi_m_valid : out STD_LOGIC;   '           axi_m_last  : out STD_LOGIC;   '           axi_m_ready : in  STD_LOGIC;       <           axi_s_data  : in  STD_LOGIC_VECTOR (7  downto 0);   '           axi_s_valid : in  STD_LOGIC;   '           axi_s_last  : in  STD_LOGIC;   '           axi_s_ready : out STD_LOGIC;�      	   Q      <           axi_m_data  : out STD_LOGIC_VECTOR (7  downto 0);5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                V       ^
f   1 �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      "   --s_ready           <= emi(13);�   L   N   Q         emo(12)           <= s_last;�   K   M   Q          emo(11)           <= s_valid;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);�   H   J   Q          emo(10)           <= m_ready;�   G   I   Q         m_last            <= emi(9);�   F   H   Q      "   --`m_valid           <= emi(8);�   E   G   Q      (   m_data            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q                     s_ready <= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      &                  last_s_ready <= '1';�   8   :   Q      &                  s_ready      <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q                     m_valid <= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      &                  last_m_valid <= '1';�   #   %   Q      &                  m_valid      <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      8           emo     : out STD_LOGIC_VECTOR (31 downto 0);�         Q      8           emi     : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �                7           leds    : out STD_LOGIC_VECTOR (3 downto 0);�                (           axi_s_tlast  : in  STD_LOGIC;�                "           clk     : in STD_LOGIC;�                (           axi_s_tvalid : in  STD_LOGIC;�                =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
             (           axi_m_tready : in  STD_LOGIC;�   	             (           axi_m_tlast  : out STD_LOGIC;�                (           axi_s_tready : out STD_LOGIC;�      	          =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�                #           rst     : in STD_LOGIC);5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                                                V       ^'     �   #   %   Q      &                  m_valid      <= '1';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                                                V       ^'     �   #   %   Q      &                  m_valid      <= '1';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                                                V       ^'     �   #   %   Q      1                  m_axis_tvalidvalid      <= '1';5�_�  �  �  �      �   $        ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^'#     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      "   --s_ready           <= emi(13);�   L   N   Q         emo(12)           <= s_last;�   K   M   Q          emo(11)           <= s_valid;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);�   H   J   Q          emo(10)           <= m_ready;�   G   I   Q         m_last            <= emi(9);�   F   H   Q      "   --`m_valid           <= emi(8);�   E   G   Q      (   m_data            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q                     s_ready <= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      &                  last_s_ready <= '1';�   8   :   Q      &                  s_ready      <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q                     m_valid <= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   #   %          &                  m_axis_tvalid<= '1';�   $   &          &                  last_m_valid <= '1';5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^''     �   '   )   Q                     m_valid <= '0';5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^'*     �   '   )   Q      )               m_axis_tvalidvalid <= '0';5�_�  �  �          �   (        ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^',     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      "   --s_ready           <= emi(13);�   L   N   Q         emo(12)           <= s_last;�   K   M   Q          emo(11)           <= s_valid;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);�   H   J   Q          emo(10)           <= m_ready;�   G   I   Q         m_last            <= emi(9);�   F   H   Q      "   --`m_valid           <= emi(8);�   E   G   Q      (   m_data            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q                     s_ready <= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      &                  last_s_ready <= '1';�   8   :   Q      &                  s_ready      <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   '   )          #               m_axis_tvalid<= '0';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^'3     �   8   :   Q      &                  s_ready      <= '1';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^'6     �   8   :   Q      1                  s_axis_treadyready      <= '1';5�_�  �  �          �   9        ����                                                                                                                                                                                                                                                                                                                            9          :          V       ^'8     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      "   --s_ready           <= emi(13);�   L   N   Q         emo(12)           <= s_last;�   K   M   Q          emo(11)           <= s_valid;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);�   H   J   Q          emo(10)           <= m_ready;�   G   I   Q         m_last            <= emi(9);�   F   H   Q      "   --`m_valid           <= emi(8);�   E   G   Q      (   m_data            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q                     s_ready <= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      '                  last_s_ready  <= '1';�   8   :   Q      '                  s_axis_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   8   :          &                  s_axis_tready<= '1';�   9   ;          &                  last_s_ready <= '1';5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            9          :          V       ^'=     �   <   >   Q                     s_ready <= '0';5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            9          :          V       ^'?     �   <   >   Q      )               s_axis_treadyready <= '0';5�_�  �  �          �   =        ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'A     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      "   --s_ready           <= emi(13);�   L   N   Q         emo(12)           <= s_last;�   K   M   Q          emo(11)           <= s_valid;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);�   H   J   Q          emo(10)           <= m_ready;�   G   I   Q         m_last            <= emi(9);�   F   H   Q      "   --`m_valid           <= emi(8);�   E   G   Q      (   m_data            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      #               s_axis_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      '                  last_s_ready  <= '1';�   8   :   Q      '                  s_axis_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   <   >          #               s_axis_tready<= '0';5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'H     �   F   H   Q      "   --`m_valid           <= emi(8);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'H     �   F   H   Q      !   -`m_valid           <= emi(8);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'I     �   F   H   Q          `m_valid           <= emi(8);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'J     �   F   H   Q         m_valid           <= emi(8);5�_�  �  �          �   N   "    ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'M     �   M   O   Q      "   --s_ready           <= emi(13);5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'O     �   M   O   Q      %   --s_ready           <= emi(13); --5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                            =          =          V       ^'O     �   M   O   Q      $   -s_ready           <= emi(13); --5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^'T     �   F   I   Q      "   m_valid           <= emi(8); --      m_last            <= emi(9);�   E   G   Q      (   m_data            <= emi(7 downto 0);5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^'`     �   K   N   Q          emo(11)           <= s_valid;      emo(12)           <= s_last;�   J   L   Q      +   emo(7   downto 0) <= s_data(7 downto 0);5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^'d     �   H   J   Q          emo(10)           <= m_ready;5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^'s     �   M   O   Q      #   s_ready           <= emi(13); --5�_�  �  �          �   K        ����                                                                                                                                                                                                                                                                                                                            N   
       K   
       V   
    ^'{     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      #   s_axi_tready      <= emi(13); --�   L   N   Q      $   emo(12)           <= s_axi_tlast;�   K   M   Q      %   emo(11)           <= s_axi_tvalid;�   J   L   Q      0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);�   H   J   Q      %   emo(10)           <= m_axi_tready;�   G   I   Q      $   m_axi_tlast            <= emi(9);�   F   H   Q      '   m_axi_tvalid           <= emi(8); --�   E   G   Q      -   m_axi_tdata            <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      #               s_axis_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      '                  last_s_ready  <= '1';�   8   :   Q      '                  s_axis_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   J   L          0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);�   M   O          (   s_axi_tready           <= emi(13); --�   L   N          $   emo(12)           <= s_axi_tlast;�   K   M          %   emo(11)           <= s_axi_tvalid;5�_�  �  �          �   F        ����                                                                                                                                                                                                                                                                                                                            I           F           V        ^'|     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      #   s_axi_tready      <= emi(13); --�   L   N   Q      $   emo(12)           <= s_axi_tlast;�   K   M   Q      %   emo(11)           <= s_axi_tvalid;�   J   L   Q      0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);�   H   J   Q          emo(10)      <= m_axi_tready;�   G   I   Q         m_axi_tlast  <= emi(9);�   F   H   Q         m_axi_tvalid <= emi(8); --�   E   G   Q      #   m_axi_tdata  <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      #               s_axis_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      '                  last_s_ready  <= '1';�   8   :   Q      '                  s_axis_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   E   G          -   m_axi_tdata            <= emi(7 downto 0);�   H   J          %   emo(10)           <= m_axi_tready;�   G   I          $   m_axi_tlast            <= emi(9);�   F   H          '   m_axi_tvalid           <= emi(8); --5�_�  �  �          �   F        ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^'�     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      #   s_axi_tready      <= emi(13); --�   L   N   Q      $   emo(12)           <= s_axi_tlast;�   K   M   Q      %   emo(11)           <= s_axi_tvalid;�   J   L   Q      0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);�   H   J   Q      %   emo(10)           <= m_axi_tready;�   G   I   Q         m_axi_tlast       <= emi(9);�   F   H   Q      "   m_axi_tvalid      <= emi(8); --�   E   G   Q      (   m_axi_tdata       <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      #               s_axis_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      '                  last_s_ready  <= '1';�   8   :   Q      '                  s_axis_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      #               m_axis_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      '                  m_axis_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   E   G          #   m_axi_tdata  <= emi(7 downto 0);�   M   O          #   s_axi_tready      <= emi(13); --�   L   N          $   emo(12)           <= s_axi_tlast;�   K   M          %   emo(11)           <= s_axi_tvalid;�   O   Q          +   leds              <= emi(17  downto 14);�   H   J              emo(10)      <= m_axi_tready;�   G   I             m_axi_tlast  <= emi(9);�   F   H             m_axi_tvalid <= emi(8); --�   J   L          0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^'�     �   F   H   Q      "   m_axi_tvalid      <= emi(8); --5�_�  �  �          �   N       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^'�   2 �   M   O   Q      #   s_axi_tready      <= emi(13); --5�_�  �  �          �   (       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^(     �   '   )   Q      #               m_axis_tvalid<= '0';5�_�  �  �  �      �   (       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^(     �   '   )   Q      '               axi_m_axis_tvalid<= '0';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^(#     �   #   %   Q      '                  m_axis_tvalid <= '1';5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^((     �   #   %   Q      +                  axi_m_axis_tvalid <= '1';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^(3     �   8   :   Q      '                  s_axis_tready <= '1';5�_�  �  �          �   9       ����                                                                                                                                                                                                                                                                                                                            9          9          v       ^(7     �   8   :   Q      +                  axi_s_axis_tready <= '1';5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            9          9          v       ^(:     �   <   >   Q      #               s_axis_tready<= '0';5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                            =          =          v       ^(=     �   <   >   Q      '               axi+s_axis_tready<= '0';5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(C     �   F   I   Q      $   --m_axi_tvalid      <= emi(8); --      m_axi_tlast       <= emi(9);�   E   G   Q      (   m_axi_tdata       <= emi(7 downto 0);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(I     �   F   H   Q      (   axi_--m_axi_tvalid      <= emi(8); --5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(J     �   F   H   Q      '   axi_-m_axi_tvalid      <= emi(8); --5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(P     �   E   I   Q      ,   axi_m_axi_tdata       <= emi(7 downto 0);   &   axi_-_axi_tvalid      <= emi(8); --   #   axi_m_axi_tlast       <= emi(9);5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(S     �   F   H   Q      "   axi_-_tvalid      <= emi(8); --5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(U     �   F   H   Q      "   axi_m_tvalid      <= emi(8); --5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            F          H                 ^(Y     �   H   J   Q      %   emo(10)           <= m_axi_tready;5�_�  �             �   I       ����                                                                                                                                                                                                                                                                                                                            I          I           v        ^(^     �   H   J   Q      )   emo(10)           <= axi_m_axi_tready;5�_�  �                K       ����                                                                                                                                                                                                                                                                                                                            K          M                 ^(b     �   J   N   Q      0   emo(7   downto 0) <= s_axi_tdata(7 downto 0);   %   emo(11)           <= s_axi_tvalid;   $   emo(12)           <= s_axi_tlast;5�_�                  K       ����                                                                                                                                                                                                                                                                                                                            K          M                 ^(b     �   J   O   Q      ,   emo(7   downto 0) <= s_tdata(7 downto 0);   !   emo(11)           <= s_tvalid;       emo(12)           <= s_tlast;   %   --s_axi_tready      <= emi(13); --�   K   L   Q    5�_�                 N       ����                                                                                                                                                                                                                                                                                                                            K          M                 ^(i     �   M   O   Q      %   --s_axi_tready      <= emi(13); --5�_�               9        ����                                                                                                                                                                                                                                                                                                                            9          :          V       ^(z     �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      '   --s_axi_s_tready      <= emi(13); --�   L   N   Q      $   emo(12)           <= axi_s_tlast;�   K   M   Q      %   emo(11)           <= axi_s_tvalid;�   J   L   Q      0   emo(7   downto 0) <= axi_s_tdata(7 downto 0);�   H   J   Q      %   emo(10)           <= axi_m_tready;�   G   I   Q         axi_m_tlast       <= emi(9);�   F   H   Q      $   --axi_m_tvalid      <= emi(8); --�   E   G   Q      (   axi_m_tdata       <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      "               axi+s_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      &                  last_s_ready <= '1';�   8   :   Q      &                  axi_s_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      "               axi_m_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      '                  last_m_valid  <= '1';�   #   %   Q      &                  axi_m_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   8   :          &                  axi_s_tready <= '1';�   9   ;          '                  last_s_ready  <= '1';5�_�                 $        ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^(~   3 �   O   Q   Q      +   leds              <= emi(17  downto 14);�   M   O   Q      '   --s_axi_s_tready      <= emi(13); --�   L   N   Q      $   emo(12)           <= axi_s_tlast;�   K   M   Q      %   emo(11)           <= axi_s_tvalid;�   J   L   Q      0   emo(7   downto 0) <= axi_s_tdata(7 downto 0);�   H   J   Q      %   emo(10)           <= axi_m_tready;�   G   I   Q         axi_m_tlast       <= emi(9);�   F   H   Q      $   --axi_m_tvalid      <= emi(8); --�   E   G   Q      (   axi_m_tdata       <= emi(7 downto 0);�   C   E   Q         end process s_one_shot;�   B   D   Q            end if;�   A   C   Q               end if;�   @   B   Q                  end if;�   ?   A   Q                     end if;�   >   @   Q      &                  last_s_ready <= '0';�   =   ?   Q      #               if(emi(13)='0') then�   <   >   Q      "               axi+s_tready<= '0';�   ;   =   Q                  else �   :   <   Q                     end if;�   9   ;   Q      &                  last_s_ready <= '1';�   8   :   Q      &                  axi_s_tready <= '1';�   7   9   Q      #               if(emi(13)='1') then�   6   8   Q      (            if (last_s_ready = '0') then�   5   7   Q               else �   4   6   Q                  last_s_ready <='0';�   3   5   Q               if rst='0' then�   2   4   Q            if rising_edge(clk) then�   1   3   Q         begin�   0   2   Q         s_one_shot:process(clk) is�   .   0   Q         end process m_one_shot;�   -   /   Q            end if;�   ,   .   Q               end if;�   +   -   Q                  end if;�   *   ,   Q                     end if;�   )   +   Q      &                  last_m_valid <= '0';�   (   *   Q      "               if(emi(8)='0') then�   '   )   Q      "               axi_m_tvalid<= '0';�   &   (   Q                  else �   %   '   Q                     end if;�   $   &   Q      &                  last_m_valid <= '1';�   #   %   Q      &                  axi_m_tvalid <= '1';�   "   $   Q      "               if(emi(8)='1') then�   !   #   Q      (            if (last_m_valid = '0') then�       "   Q               else �      !   Q                  last_m_valid <='0';�          Q               if rst='0' then�         Q            if rising_edge(clk) then�         Q         begin�         Q         m_one_shot:process(clk) is�         Q      +      signal last_s_ready: STD_LOGIC :='0';�         Q      +      signal last_m_valid: STD_LOGIC :='0';�         Q      )           rst          : in  STD_LOGIC);�         Q      =           leds         : out STD_LOGIC_VECTOR (3  downto 0);�         Q      (           clk          : in  STD_LOGIC;�         Q      (           axi_s_tready : out STD_LOGIC;�         Q      (           axi_s_tlast  : in  STD_LOGIC;�         Q      (           axi_s_tvalid : in  STD_LOGIC;�         Q      =           axi_s_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�   
      Q      (           axi_m_tready : in  STD_LOGIC;�   	      Q      (           axi_m_tlast  : out STD_LOGIC;�      
   Q      (           axi_m_tvalid : out STD_LOGIC;�      	   Q      =           axi_m_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�         Q      =           emo          : out STD_LOGIC_VECTOR (31 downto 0);�         Q      =           emi          : in  STD_LOGIC_VECTOR (31 downto 0);�         Q          Port(  �   #   %          &                  axi_m_tvalid <= '1';�   $   &          '                  last_m_valid  <= '1';5�_�                 =       ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^(�     �   <   >   Q      "               axi+s_tready<= '0';5�_�                   =       ����                                                                                                                                                                                                                                                                                                                            $           %           V        ^(�   4 �   <   >   Q      "               axi+s_tready<= '0';5�_�                 9        ����                                                                                                                                                                                                                                                                                                                            9          :          V       ^(u     �   8   ;   Q      &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   'eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �  �      �  �   (       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^(     �   '   )   Q                     axi_m<= '0';5�_�  �              �   (       ����                                                                                                                                                                                                                                                                                                                            F           Q           V        ^(     �   '   )   Q                     axi_uum<= '0';5�_�  �          �  �   $        ����                                                                                                                                                                                                                                                                                                                            $          %          V       ^'      �   #   &   Q      &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �          �  �   9       ����                                                                                                                                                                                                                                                                                                                         :          B          V       ^�U     �   8   :   U                  last_s_ready <=0'';5�_�  �          �  �   8   	    ����                                                                                                                                                                                                                                                                                                                         #   	       %   	       V   	    ^��     �   7   :   W      +         if rst='0' then last_m_valid <=0';5�_�  �  �      �  �   $       ����                                                                                                                                                                                                                                                                                                                                             V       ^��     �   $   %   R    �   #   $   R      +      signal last_s_ready: STD_LOGIC :='0';   begin5�_�  �              �   $       ����                                                                                                                                                                                                                                                                                                                                             V       ^��     �   #   %   T      1            signal last_s_ready: STD_LOGIC :='0';5�_�  �          �  �      
    ����                                                                                                                                                                                                                                                                                                                                               V        ^�G     �         N            �         O            kllllll5�_�  K          M  L   $       ����                                                                                                                                                                                                                                                                                                                         "          "          v       ^��     �   $   %   7    �   #   %   7      "        lrising_edge(emi(8)) then 5�_�  $          &  %          ����                                                                0                                                                                                                                             0                                                                                                          2           2          V   ,    ^�;     �         5      <           s_clk   : out STD_LOGIC; s_clk   : out STD_LOGIC;5�_�            	            ����                                                                                                                                                                                                                                                                                                                           )   %       )   (       v   (    ^�^     �         )          �         *          j5�_�   �       �   �   �   )       ����                                                                                                                                                    ,                                                                                                                                                                                          V   ,    ^�     �   (   )   ,       5�_�   �           �   �   )       ����                                                                                                                                                    ,                                                                                                                                                                                          V   ,    ^�     �   (   )   ,         �   (   *   -         h5�_�   e           g   f           ����                                                                                                                                                                                                                                                                                                                                         
       v   
    ^��     �      !   #         s<S-F11>emo(10)  <= m_ready;5�_�   1   3       4   2          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^~�     �   
            $           m_clk   : in   STD_LOGIC;5�_�   2               3          ����                                                                                                                                                                                                                                                                                                                            
   $          $          $    ^~�     �   
            %           m_clk   : in    STD_LOGIC;5�_�   )           +   *          ����                                                                                                                                                                                                                                                                                                                                                V       ^}7     �                   <= emio(8);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^|0     �               B    Port( emo :                in  STD_LOGIC_VECTOR (15 downto 0);5��