Vim�UnDo� �~�,X%Y�J=�/2�L�6�.9t[�0��   >                                   ^�    _�                              ����                                                                                                                                                                                                                                                                                                                                                             ^�    �                'architecture Behavioral of join_8to2 is�                end join_8to2;�                entity join_8to2 is5��