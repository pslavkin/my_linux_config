Vim�UnDo� �����Uv��|�a@���Rj��ܗ�3&&   @                0      0  0  0    ^N�    _�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ^
p    �               *           rst           : in  STD_LOGIC);�               "           clk     : in STD_LOGIC;�               )           s_axis_tready : out STD_LOGIC;�               )           s_axis_tlast  : in  STD_LOGIC;�               )           s_axis_tvalid : in  STD_LOGIC;�   
            =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
         )           m_axis_tready : in  STD_LOGIC;�      	         )           m_axis_tlast  : out STD_LOGIC;�               )           m_axis_tvalid : out STD_LOGIC;�               >           m_axis_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�                   Port(  �                #           rst     : in STD_LOGIC);�                )           s_axis_tready : out STD_LOGIC;�                )           s_axis_tlast  : in  STD_LOGIC;�   
             >           s_axis_tdata  : in  STD_LOGIC_VECTOR (7  downto 0);�      	          )           m_axis_tlast  : out STD_LOGIC;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �                  �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�    �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �                     �             5�_�                          ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �               	         �             5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �                        if rst = '1'5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �                        if rst = '0'5�_�   	              
      
    ����                                                                                                                                                                                                                                                                                                                                                  V        ^J     �         !                  �              5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                  V        ^Z     �         #         �         "    5�_�                      +    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         #      +   signal state:STD_LOGIC_VECTOR (3 downto 5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         #      <   signal state:STD_LOGIC_VECTOR (3 downto 0):= others=>'0')5�_�                       =    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         #      =   signal state:STD_LOGIC_VECTOR (3 downto 0):= (others=>'0')5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       "   #         end process shift_reg;�          #               end if;�         #               else�         #                  bitCounter:=0;�         #               if rst = '0' then�         #            if rising_edge(clk) then�         #         begin�         #         shift_reg:process (clk) is�         #      @   signal state:STD_LOGIC_VECTOR ( 3 downto 0 ):= (others=>'0');�         #      *           rst           : in  STD_LOGIC);�         #      )           clk           : in  STD_LOGIC;�         #      )           s_axis_tready : out STD_LOGIC;�         #      )           s_axis_tlast  : in  STD_LOGIC;�         #      )           s_axis_tvalid : in  STD_LOGIC;�   
      #      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   #      )           m_axis_tready : in  STD_LOGIC;�      	   #      )           m_axis_tlast  : out STD_LOGIC;�         #      )           m_axis_tvalid : out STD_LOGIC;�         #      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         #          Port(  �                >   signal state:STD_LOGIC_VECTOR (3 downto 0):= (others=>'0');5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         #       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         #       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �                 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         "    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         #                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^U     �         #      #            m_axis_tdata(0)        5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^V     �         #                  m_axis_tdata(0)5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^X     �         #                  m_axis_tdata(0)l5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^_     �         #                  m_axis_tdata(0);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �          $                  �          #    5�_�                       &    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �      !   $    5�_�                             ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �                  5�_�                       	    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �         %                  �         $    5�_�                         !    ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       "   &                  �       "   %    5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                	          	       V   	    ^�     �   #   %   &         end process shift_reg;�   !   #   &               end if;�       "   &               end if;�      !   &      ,            bitCounter      := bitCounter+1;�          &      8            m_axis_tdata(0) <= s_axis_tdata(bitCounter);�         &      "            if bitCounter < 8 then�         &               else�         &                  bitCounter:=0;�         &               if rst = '0' then�         &            if rising_edge(clk) then�         &         begin�         &         shift_reg:process (clk) is�         &      @   signal state:STD_LOGIC_VECTOR ( 3 downto 0 ):= (others=>'0');�         &      *           rst           : in  STD_LOGIC);�         &      )           clk           : in  STD_LOGIC;�         &      )           s_axis_tready : out STD_LOGIC;�         &      )           s_axis_tlast  : in  STD_LOGIC;�         &      )           s_axis_tvalid : in  STD_LOGIC;�   
      &      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   &      )           m_axis_tready : in  STD_LOGIC;�      	   &      )           m_axis_tlast  : out STD_LOGIC;�         &      )           m_axis_tvalid : out STD_LOGIC;�         &      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         &          Port(  �                 8            m_axis_tdata(0) <= s_axis_tdata(bitCounter);�      !          '            bitCounter := bitCounter+1;5�_�       "           !   !        ����                                                                                                                                                                                                                                                                                                                                	          	       V   	    ^�     �       "   &               end if;5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �      !          ,            bitCounter      := bitCounter+1;�                 8            m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   "   $           #   #        ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �   "   $   &    �   #   $   &    5�_�   #   %           $   #       ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �   "   $                   end if;5�_�   $   &           %   $        ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �   #   $           5�_�   %   '           &   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �       "   &                  end if;5�_�   &   (           '   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �       #   &                  e5�_�   '   )           (   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �   !   #   '                     m_axis_tvalid5�_�   (   *           )           ����                                                                                                                                                                                                                                                                                                                                                 V       ^�     �         (         �         '    5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                            !                     V       ^     �         (         type state5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                            !                     V       ^     �         (         type shiftSstate5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                            !                     V       ^     �         (         type shiftState5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                v       ^?     �         (      @   signal state:STD_LOGIC_VECTOR ( 3 downto 0 ):= (others=>'0');5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                         (       v   (    ^E     �         (      :   signal state:shiftState ( 3 downto 0 ):= (others=>'0');5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^H     �         (      ,   signal state:shiftState := (others=>'0');5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^X     �         (    �         (    5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^Y     �         )                  bitCounter:=0;5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^^     �         )                  state:=0;5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^`     �         )                  state<=0;5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^a     �         )                  state<=idle0;5�_�   4   7           5           ����                                                                                                                                                                                                                                                                                                                                                V       ^e     �   &   (   )         end process shift_reg;�   %   '   )            end if;�   $   &   )               end if;�   #   %   )      !               m_axis_tvalid <=0;�   "   $   )                  else�   !   #   )      /               bitCounter      := bitCounter+1;�       "   )      ;               m_axis_tdata(0) <= s_axis_tdata(bitCounter);�      !   )      "            if bitCounter < 8 then�          )               else�         )                  bitCounter := 0;�         )                  state      <= idle;�         )               if rst = '0' then�         )            if rising_edge(clk) then�         )         begin�         )         shift_reg:process (clk) is�         )      #   signal state:shiftState := idle;�         )      '   type shiftState is (idle, shifting);�         )      *           rst           : in  STD_LOGIC);�         )      )           clk           : in  STD_LOGIC;�         )      )           s_axis_tready : out STD_LOGIC;�         )      )           s_axis_tlast  : in  STD_LOGIC;�         )      )           s_axis_tvalid : in  STD_LOGIC;�   
      )      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   )      )           m_axis_tready : in  STD_LOGIC;�      	   )      )           m_axis_tlast  : out STD_LOGIC;�         )      )           m_axis_tvalid : out STD_LOGIC;�         )      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         )          Port(  �                            state<=idle;�                            bitCounter:=0;5�_�   5   8   6       7           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �      "   *                  �      !   )    5�_�   7   9           8   !       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       "   +    5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �      !   ,    5�_�   9   ;           :   !       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       "   -    �   !   "   -    5�_�   :   <           ;            ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �                  5�_�   ;   =           <   !       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       !                      case state is5�_�   <   >           =   !        ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       !           5�_�   =   ?           >   !       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �       "   +    �   !   "   +    5�_�   >   @           ?   "       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �   !   #   ,                     when idle =>5�_�   ?   A           @   "       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �   "   $   -                        �   "   $   ,    5�_�   @   B           A   $        ����                                                                                                                                                                                                                                                                                                                            $          )          V       ^     �   #   $          "            if bitCounter < 8 then   ;               m_axis_tdata(0) <= s_axis_tdata(bitCounter);   /               bitCounter      := bitCounter+1;               else   !               m_axis_tvalid <=0;            end if;5�_�   A   C           B   #       ����                                                                                                                                                                                                                                                                                                                            $          $          V       ^     �   "   )   '    �   #   $   '    5�_�   B   D           C   #        ����                                                                                                                                                                                                                                                                                                                            #          '          V       ^     �   &   (          !               m_axis_tvalid <=0;�   %   '                      else�   $   &          /               bitCounter      := bitCounter+1;�   #   %          ;               m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   "   $          "            if bitCounter < 8 then5�_�   C   E           D   "       ����                                                                                                                                                                                                                                                                                                                            #          '          V       ^     �   !   #   -    �   "   #   -    5�_�   D   F           E   "       ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^     �   !   #   .      (                  if bitCounter < 8 then5�_�   E   G           F   "       ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^+     �   !   #   .      +                  if m_axis_tvalid < 8 then5�_�   F   H           G   "   #    ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^/     �   !   #   .      +                  if m_axis_tready < 8 then5�_�   G   I           H   "   $    ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^/     �   !   #   .      ,                  if m_axis_tready =< 8 then5�_�   H   J           I   "   %    ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^1     �   !   #   .      +                  if m_axis_tready = 8 then5�_�   I   K           J   "   (    ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^2     �   !   #   .      .                  if m_axis_tready = '1'8 then5�_�   J   L           K   "   (    ����                                                                                                                                                                                                                                                                                                                            $          (          V       ^<     �   "   $   .    5�_�   K   M           L   #        ����                                                                                                                                                                                                                                                                                                                            %          )          V       ^@     �   "   $   /    �   #   $   /    5�_�   L   N           M   #   %    ����                                                                                                                                                                                                                                                                                                                            &          *          V       ^B     �   "   $   0      '                     m_axis_tvalid <=0;5�_�   M   O           N   $        ����                                                                                                                                                                                                                                                                                                                            &          *          V       ^j     �   #   %   0    �   $   %   0    5�_�   N   P           O   #        ����                                                                                                                                                                                                                                                                                                                            #          $          V       ^�     �   .   0   1         end process shift_reg;�   -   /   1            end if;�   ,   .   1                  end case;�   +   -   1               end if;�   *   ,   1      '                     m_axis_tvalid <=0;�   )   +   1                        else�   (   *   1      5                     bitCounter      := bitCounter+1;�   '   )   1      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   &   (   1      (                  if bitCounter < 8 then�   %   '   1                     when shifting =>�   #   %   1      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   "   $   1      *                     m_axis_tvalid   <= 1;�   !   #   1      -                  if m_axis_tready = '1' then�       "   1                     when idle =>�      !   1                  case state is�          1               else�         1                  bitCounter := 0;�         1                  state      <= idle;�         1               if rst = '0' then�         1            if rising_edge(clk) then�         1         begin�         1         shift_reg:process (clk) is�         1      #   signal state:shiftState := idle;�         1      '   type shiftState is (idle, shifting);�         1      *           rst           : in  STD_LOGIC);�         1      )           clk           : in  STD_LOGIC;�         1      )           s_axis_tready : out STD_LOGIC;�         1      )           s_axis_tlast  : in  STD_LOGIC;�         1      )           s_axis_tvalid : in  STD_LOGIC;�   
      1      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   1      )           m_axis_tready : in  STD_LOGIC;�      	   1      )           m_axis_tlast  : out STD_LOGIC;�         1      )           m_axis_tvalid : out STD_LOGIC;�         1      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         1          Port(  �   "   $          '                     m_axis_tvalid <=1;�   #   %          A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   O   Q           P   %        ����                                                                                                                                                                                                                                                                                                                            #          $          V       ^�     �   $   &   1    �   %   &   1    5�_�   P   R           Q   %       ����                                                                                                                                                                                                                                                                                                                            #          $          V       ^�     �   $   &   2                  state      <= idle;5�_�   Q   S           R   %       ����                                                                                                                                                                                                                                                                                                                            #          $          V       ^�     �   $   &   2      (                     state      <= idle;5�_�   R   T           S   %       ����                                                                                                                                                                                                                                                                                                                            #          $          V       ^�     �   $   &   2      #                     state <= idle;5�_�   S   U           T   #        ����                                                                                                                                                                                                                                                                                                                            %   %       #   %       V   %    ^�     �   /   1   2         end process shift_reg;�   .   0   2            end if;�   -   /   2                  end case;�   ,   .   2               end if;�   +   -   2      '                     m_axis_tvalid <=0;�   *   ,   2                        else�   )   +   2      5                     bitCounter      := bitCounter+1;�   (   *   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   '   )   2      (                  if bitCounter < 8 then�   &   (   2                     when shifting =>�   $   &   2      1                     state           <= shifting;�   #   %   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   "   $   2      *                     m_axis_tvalid   <= 1;�   !   #   2      -                  if m_axis_tready = '1' then�       "   2                     when idle =>�      !   2                  case state is�          2               else�         2                  bitCounter := 0;�         2                  state      <= idle;�         2               if rst = '0' then�         2            if rising_edge(clk) then�         2         begin�         2         shift_reg:process (clk) is�         2      #   signal state:shiftState := idle;�         2      '   type shiftState is (idle, shifting);�         2      *           rst           : in  STD_LOGIC);�         2      )           clk           : in  STD_LOGIC;�         2      )           s_axis_tready : out STD_LOGIC;�         2      )           s_axis_tlast  : in  STD_LOGIC;�         2      )           s_axis_tvalid : in  STD_LOGIC;�   
      2      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   2      )           m_axis_tready : in  STD_LOGIC;�      	   2      )           m_axis_tlast  : out STD_LOGIC;�         2      )           m_axis_tvalid : out STD_LOGIC;�         2      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         2          Port(  �   "   $          *                     m_axis_tvalid   <= 1;�   $   &          '                     state <= shifting;�   #   %          A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   T   V           U   %        ����                                                                                                                                                                                                                                                                                                                            %   %       #   %       V   %    ^�     �   %   '   3                           �   %   '   2    5�_�   U   W           V   '        ����                                                                                                                                                                                                                                                                                                                            %   %       #   %       V   %    ^�     �   &   '           5�_�   V   X           W   &       ����                                                                                                                                                                                                                                                                                                                            %   %       #   %       V   %    ^�     �   %   '   2    �   &   '   2    5�_�   W   Y           X   &       ����                                                                                                                                                                                                                                                                                                                            %   %       #   %       V   %    ^�     �   %   '                      bitCounter := 0;5�_�   X   Z           Y   #        ����                                                                                                                                                                                                                                                                                                                            &          #          V       ^�     �   0   2   3         end process shift_reg;�   /   1   3            end if;�   .   0   3                  end case;�   -   /   3               end if;�   ,   .   3      '                     m_axis_tvalid <=0;�   +   -   3                        else�   *   ,   3      5                     bitCounter      := bitCounter+1;�   )   +   3      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   (   *   3      (                  if bitCounter < 8 then�   '   )   3                     when shifting =>�   &   (   3                        end if;�   %   '   3      *                     bitCounter      := 0;�   $   &   3      1                     state           <= shifting;�   #   %   3      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   "   $   3      *                     m_axis_tvalid   <= 1;�   !   #   3      -                  if m_axis_tready = '1' then�       "   3                     when idle =>�      !   3                  case state is�          3               else�         3                  bitCounter := 0;�         3                  state      <= idle;�         3               if rst = '0' then�         3            if rising_edge(clk) then�         3         begin�         3         shift_reg:process (clk) is�         3      #   signal state:shiftState := idle;�         3      '   type shiftState is (idle, shifting);�         3      *           rst           : in  STD_LOGIC);�         3      )           clk           : in  STD_LOGIC;�         3      )           s_axis_tready : out STD_LOGIC;�         3      )           s_axis_tlast  : in  STD_LOGIC;�         3      )           s_axis_tvalid : in  STD_LOGIC;�   
      3      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   3      )           m_axis_tready : in  STD_LOGIC;�      	   3      )           m_axis_tlast  : out STD_LOGIC;�         3      )           m_axis_tvalid : out STD_LOGIC;�         3      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         3          Port(  �   "   $          *                     m_axis_tvalid   <= 1;�   %   '          %                     bitCounter := 0;�   $   &          1                     state           <= shifting;�   #   %          A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   Y   [           Z           ����                                                                                                                                                                                                                                                                                                                            &          #          V       ^�     �                            bitCounter := 0;5�_�   Z   \           [           ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �      !   2                     when idle =>5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2                  state      <= idle;5�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2      '   type shiftState is (idle, shifting);5�_�   ]   _           ^          ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2      #   signal state:shiftState := idle;5�_�   ^   `           _           ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2      &            state      <= waitinReady;5�_�   _   a           `      $    ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2      *   signal state:shiftState := waitinReady;5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^�     �         2      .   type shiftState is (waitinReady, shifting);5�_�   a   c           b           ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^     �      !   2      "               when waitinReady =>5�_�   b   d           c   (   "    ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^     �   '   )   2      (                  if bitCounter < 8 then5�_�   c   e           d   (   "    ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^     �   '   )   2      (                  if bitCounter < 7 then5�_�   d   f           e   (   "    ����                                                                                                                                                                                                                                                                                                                            %          "          V       ^(     �   '   )   2      (                  if bitCounter < 8 then5�_�   e   g           f   "        ����                                                                                                                                                                                                                                                                                                                            "   "       "   "       V   "    ^D     �   !   "          *                     m_axis_tvalid   <= 1;5�_�   f   h           g   '       ����                                                                                                                                                                                                                                                                                                                            "   "       "   "       V   "    ^L     �   &   (   1    �   '   (   1    5�_�   g   i           h   (   "    ����                                                                                                                                                                                                                                                                                                                            "   "       "   "       V   "    ^N     �   '   )   2      (                  if bitCounter < 7 then5�_�   h   j           i   '        ����                                                                                                                                                                                                                                                                                                                            '   "       '   "       V   "    ^t     �   &   '          *                     m_axis_tvalid   <= 1;5�_�   i   k           j   (       ����                                                                                                                                                                                                                                                                                                                            '   "       '   "       V   "    ^u     �   '   )   1    �   (   )   1    5�_�   j   l           k   "       ����                                                                                                                                                                                                                                                                                                                            '   "       '   "       V   "    ^�     �   !   "          A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   k   m           l   )       ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^�     �   )   +   2                           �   )   +   1    5�_�   l   n           m   *       ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^     �   )   *          '                     if(bitCounter = 8)5�_�   m   o           n   ,       ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^     �   +   -   1    �   ,   -   1    5�_�   n   p           o   ,   (    ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^      �   +   -   2      1                     state           <= shifting;5�_�   o   q           p   ,   3    ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^#     �   ,   .   3                           �   ,   .   2    5�_�   p   r           q   .   	    ����                                                                                                                                                                                                                                                                                                                            &   "       &   "       V   "    ^-     �   -   .                   end if;5�_�   q   s           r   +        ����                                                                                                                                                                                                                                                                                                                            +          ,          V       ^2     �   /   1   2         end process shift_reg;�   .   0   2            end if;�   -   /   2                  end case;�   ,   .   2                        end if;�   +   -   2      3                     state         <= waitingReady;�   *   ,   2      (                     m_axis_tvalid <= 0;�   )   +   2                        else�   (   *   2      5                     bitCounter      := bitCounter+1;�   '   )   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   &   (   2      *                     m_axis_tvalid   <= 1;�   %   '   2      (                  if bitCounter < 8 then�   $   &   2                     when shifting =>�   #   %   2                        end if;�   "   $   2      *                     bitCounter      := 0;�   !   #   2      1                     state           <= shifting;�       "   2      -                  if m_axis_tready = '1' then�      !   2      #               when waitingReady =>�          2                  case state is�         2               else�         2      '            state      <= waitingReady;�         2               if rst = '0' then�         2            if rising_edge(clk) then�         2         begin�         2         shift_reg:process (clk) is�         2      +   signal state:shiftState := waitingReady;�         2      /   type shiftState is (waitingReady, shifting);�         2      *           rst           : in  STD_LOGIC);�         2      )           clk           : in  STD_LOGIC;�         2      )           s_axis_tready : out STD_LOGIC;�         2      )           s_axis_tlast  : in  STD_LOGIC;�         2      )           s_axis_tvalid : in  STD_LOGIC;�   
      2      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   2      )           m_axis_tready : in  STD_LOGIC;�      	   2      )           m_axis_tlast  : out STD_LOGIC;�         2      )           m_axis_tvalid : out STD_LOGIC;�         2      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         2          Port(  �   *   ,          '                     m_axis_tvalid <=0;�   +   -          5                     state           <= waitingReady;5�_�   r   t           s           ����                                                                                                                                                                                                                                                                                                                                                  V        ^8     �   /   1   2         end process shift_reg;�   .   0   2            end if;�   -   /   2                  end case;�   ,   .   2                        end if;�   +   -   2      3                     state         <= waitingReady;�   *   ,   2      (                     m_axis_tvalid <= 0;�   )   +   2                        else�   (   *   2      5                     bitCounter      := bitCounter+1;�   '   )   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   &   (   2      *                     m_axis_tvalid   <= 1;�   %   '   2      (                  if bitCounter < 8 then�   $   &   2                     when shifting =>�   #   %   2                        end if;�   "   $   2      *                     bitCounter      := 0;�   !   #   2      1                     state           <= shifting;�       "   2      -                  if m_axis_tready = '1' then�      !   2      #               when waitingReady =>�          2                  case state is�         2               else�         2      "            state <= waitingReady;�         2               if rst = '0' then�         2            if rising_edge(clk) then�         2         begin�         2         shift_reg:process (clk) is�         2      +   signal state:shiftState := waitingReady;�         2      /   type shiftState is (waitingReady, shifting);�         2      *           rst           : in  STD_LOGIC);�         2      )           clk           : in  STD_LOGIC;�         2      )           s_axis_tready : out STD_LOGIC;�         2      )           s_axis_tlast  : in  STD_LOGIC;�         2      )           s_axis_tvalid : in  STD_LOGIC;�   
      2      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   2      )           m_axis_tready : in  STD_LOGIC;�      	   2      )           m_axis_tlast  : out STD_LOGIC;�         2      )           m_axis_tvalid : out STD_LOGIC;�         2      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         2          Port(  �                '            state      <= waitingReady;5�_�   s   u           t   "        ����                                                                                                                                                                                                                                                                                                                            "           #           V        ^<     �   /   1   2         end process shift_reg;�   .   0   2            end if;�   -   /   2                  end case;�   ,   .   2                        end if;�   +   -   2      3                     state         <= waitingReady;�   *   ,   2      (                     m_axis_tvalid <= 0;�   )   +   2                        else�   (   *   2      5                     bitCounter      := bitCounter+1;�   '   )   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   &   (   2      *                     m_axis_tvalid   <= 1;�   %   '   2      (                  if bitCounter < 8 then�   $   &   2                     when shifting =>�   #   %   2                        end if;�   "   $   2      %                     bitCounter := 0;�   !   #   2      ,                     state      <= shifting;�       "   2      -                  if m_axis_tready = '1' then�      !   2      #               when waitingReady =>�          2                  case state is�         2               else�         2      "            state <= waitingReady;�         2               if rst = '0' then�         2            if rising_edge(clk) then�         2         begin�         2         shift_reg:process (clk) is�         2      +   signal state:shiftState := waitingReady;�         2      /   type shiftState is (waitingReady, shifting);�         2      *           rst           : in  STD_LOGIC);�         2      )           clk           : in  STD_LOGIC;�         2      )           s_axis_tready : out STD_LOGIC;�         2      )           s_axis_tlast  : in  STD_LOGIC;�         2      )           s_axis_tvalid : in  STD_LOGIC;�   
      2      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   2      )           m_axis_tready : in  STD_LOGIC;�      	   2      )           m_axis_tlast  : out STD_LOGIC;�         2      )           m_axis_tvalid : out STD_LOGIC;�         2      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         2          Port(  �   !   #          1                     state           <= shifting;�   "   $          *                     bitCounter      := 0;5�_�   t   v           u   +        ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�     �   *   +          (                     m_axis_tvalid <= 0;5�_�   u   w           v   !       ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�     �       "   1    �   !   "   1    5�_�   v   x           w   !       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �       "   2      (                     m_axis_tvalid <= 0;5�_�   w   y           x   !       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �       "   2      '                    m_axis_tvalid <= 0;5�_�   x   z           y   !       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �       "   2      &                   m_axis_tvalid <= 0;5�_�   y   {           z   (        ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^�     �   '   (          *                     m_axis_tvalid   <= 1;5�_�   z   |           {   ,       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^�     �   +   -   1    �   ,   -   1    5�_�   {   }           |   +        ����                                                                                                                                                                                                                                                                                                                            +          ,          V       ^�     �   /   1   2         end process shift_reg;�   .   0   2            end if;�   -   /   2                  end case;�   ,   .   2                        end if;�   +   -   2      (                     m_axis_tvalid <= 1;�   *   ,   2      3                     state         <= waitingReady;�   )   +   2                        else�   (   *   2      5                     bitCounter      := bitCounter+1;�   '   )   2      A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   &   (   2      (                  if bitCounter < 8 then�   %   '   2                     when shifting =>�   $   &   2                        end if;�   #   %   2      %                     bitCounter := 0;�   "   $   2      ,                     state      <= shifting;�   !   #   2      -                  if m_axis_tready = '1' then�       "   2      %                  m_axis_tvalid <= 0;�      !   2      #               when waitingReady =>�          2                  case state is�         2               else�         2      "            state <= waitingReady;�         2               if rst = '0' then�         2            if rising_edge(clk) then�         2         begin�         2         shift_reg:process (clk) is�         2      +   signal state:shiftState := waitingReady;�         2      /   type shiftState is (waitingReady, shifting);�         2      *           rst           : in  STD_LOGIC);�         2      )           clk           : in  STD_LOGIC;�         2      )           s_axis_tready : out STD_LOGIC;�         2      )           s_axis_tlast  : in  STD_LOGIC;�         2      )           s_axis_tvalid : in  STD_LOGIC;�   
      2      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   2      )           m_axis_tready : in  STD_LOGIC;�      	   2      )           m_axis_tlast  : out STD_LOGIC;�         2      )           m_axis_tvalid : out STD_LOGIC;�         2      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         2          Port(  �   *   ,          3                     state         <= waitingReady;�   +   -          *                     m_axis_tvalid   <= 1;5�_�   |              }          ����                                                                                                                                                                                                                                                                                                                            +          ,          V       ^e     �         2      /   type shiftState is (waitingReady, shifting);5�_�   }   �   ~                 ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ^~     �         2      +   signal state:shiftState := waitingReady;�         2    5�_�      �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        ^�     �         2      "            state <= waitingReady;�         2    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �      !   2      #               when waitingReady =>5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �       "   2      %                  m_axis_tvalid <= 0;5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �       "   2      %                  s_axis_tvalid <= 0;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �   !   #   2      -                  if m_axis_tready = '1' then5�_�   �   �   �       �   "       ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �   !   #   2      -                  if s_axis_tready = '1' then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �      !   2      %               when waitingS_Valid =>5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �      !   2      $               when waitingSValid =>5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �      !   2      $               when waitingScalid =>5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �         2      $            state <= waitingS_Valid;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �         2      #            state <= waitingSValid;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �         2      "            state <= waitingSalid;5�_�   �   �   �       �      &    ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �         2      -   signal state:shiftState := waitingS_Valid;5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    ^�     �         2      ,   signal state:shiftState := waitingSValid;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               &          &       v   &    ^�     �         2      1   type shiftState is (waitingS_Valid, shifting);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �         2      0   type shiftState is (waitingSValid, shifting);5�_�   �   �           �   +   -    ����                                                                                                                                                                                                                                                                                                                                                v       ^     �   *   ,   2      3                     state         <= waitingReady;5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                                                v       ^     �   +   -   2      (                     m_axis_tvalid <= 1;5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                                                v       ^      �   +   -   2      (                     s_axis_tvalid <= 1;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                v       ^d     �   %   '   2                     when shifting =>5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                v       ^k     �   %   '   2                     when sending =>5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                                                v       ^~     �   &   (   2    �   '   (   2    5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   &   (   3      -                  if s_axis_tvalid = '1' then5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   &   (   3      -                  if m_axis_tvalid = '1' then5�_�   �   �           �   '   #    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   *   4                           �   '   )   3    5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   (           5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   (           5�_�   �   �           �   #   #    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   "   $   3      ,                     state      <= shifting;5�_�   �   �           �   '   ,    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   )   4                           �   '   )   3    5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   (          '                     state <= shifting;5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   '   )          (                  if bitCounter < 8 then5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *          A                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   3    �   )   *   3    5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      %                  s_axis_tready <= 0;5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      +                        s_axis_tready <= 0;5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      +                        m_axis_tready <= 0;5�_�   �   �           �   )   )    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      +                        m_axis_tvalid <= 0;5�_�   �   �           �   )   )    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      +                        m_axis_tvalid <= 1;5�_�   �   �           �   )   +    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   (   *   4      ,                        m_axis_tvalid <= '1;5�_�   �   �           �   !   #    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �       "   4      %                  s_axis_tready <= 0;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �       "   4      &                  s_axis_tready <= '0;5�_�   �   �           �   $   #    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   #   %   4      %                     bitCounter := 0;5�_�   �   �           �   $   %    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   #   %   4      &                     bitCounter := '0;5�_�   �   �   �       �   )        ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^e     �   1   3   4         end process shift_reg;�   0   2   4            end if;�   /   1   4                  end case;�   .   0   4                        end if;�   -   /   4      (                     s_axis_tready <= 1;�   ,   .   4      4                     state         <= waitingSvalid;�   +   -   4                        else�   *   ,   4      5                     bitCounter      := bitCounter+1;�   )   +   4      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   (   *   4      /                        m_axis_tvalid   <= '1';�   '   )   4      +                     if bitCounter < 8 then�   &   (   4      -                  if m_axis_tready = '1' then�   %   '   4      $               when waitingMready =>�   $   &   4                        end if;�   #   %   4      '                     bitCounter := '0';�   "   $   4      1                     state      <= waitingMready;�   !   #   4      -                  if s_axis_tvalid = '1' then�       "   4      '                  s_axis_tready <= '0';�      !   4      $               when waitingSvalid =>�          4                  case state is�         4               else�         4      #            state <= waitingSvalid;�         4               if rst = '0' then�         4            if rising_edge(clk) then�         4         begin�         4         shift_reg:process (clk) is�         4      ,   signal state:shiftState := waitingSvalid;�         4      0   type shiftState is (waitingSvalid, shifting);�         4      *           rst           : in  STD_LOGIC);�         4      )           clk           : in  STD_LOGIC;�         4      )           s_axis_tready : out STD_LOGIC;�         4      )           s_axis_tlast  : in  STD_LOGIC;�         4      )           s_axis_tvalid : in  STD_LOGIC;�   
      4      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   4      )           m_axis_tready : in  STD_LOGIC;�      	   4      )           m_axis_tlast  : out STD_LOGIC;�         4      )           m_axis_tvalid : out STD_LOGIC;�         4      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         4          Port(  �   (   *          -                        m_axis_tvalid <= '1';�   )   +          D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^k     �   *   ,          5                     bitCounter      := bitCounter+1;5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^n     �   +   -                            else5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^}     �   /   1   4    �   0   1   4    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^�     �   /   1          /                        m_axis_tvalid   <= '1';5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^�     �   /   1   5      )                  m_axis_tvalid   <= '1';5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^�     �   .   0   5                        end if;5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^�     �   .   0   5                        else if;5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            )   &       *   &       V   &    ^�     �   0   2   6                           �   0   2   5    5�_�   �   �           �   0        ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^�     �   3   5   6         end process shift_reg;�   2   4   6            end if;�   1   3   6                  end case;�   0   2   6                        end if;�   /   1   6      *                     m_axis_tvalid <= '1';�   .   0   6                        else�   -   /   6      (                     s_axis_tready <= 1;�   ,   .   6      4                     state         <= waitingSvalid;�   +   -   6                           else�   *   ,   6      8                        bitCounter      := bitCounter+1;�   )   +   6      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   (   *   6      /                        m_axis_tvalid   <= '1';�   '   )   6      +                     if bitCounter < 8 then�   &   (   6      -                  if m_axis_tready = '1' then�   %   '   6      $               when waitingMready =>�   $   &   6                        end if;�   #   %   6      '                     bitCounter := '0';�   "   $   6      1                     state      <= waitingMready;�   !   #   6      -                  if s_axis_tvalid = '1' then�       "   6      '                  s_axis_tready <= '0';�      !   6      $               when waitingSvalid =>�          6                  case state is�         6               else�         6      #            state <= waitingSvalid;�         6               if rst = '0' then�         6            if rising_edge(clk) then�         6         begin�         6         shift_reg:process (clk) is�         6      ,   signal state:shiftState := waitingSvalid;�         6      0   type shiftState is (waitingSvalid, shifting);�         6      *           rst           : in  STD_LOGIC);�         6      )           clk           : in  STD_LOGIC;�         6      )           s_axis_tready : out STD_LOGIC;�         6      )           s_axis_tlast  : in  STD_LOGIC;�         6      )           s_axis_tvalid : in  STD_LOGIC;�   
      6      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   6      )           m_axis_tready : in  STD_LOGIC;�      	   6      )           m_axis_tlast  : out STD_LOGIC;�         6      )           m_axis_tvalid : out STD_LOGIC;�         6      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         6          Port(  �   /   1          ,                     m_axis_tvalid   <= '1';5�_�   �   �           �   -        ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^�     �   -   /          (                     s_axis_tready <= 1;�   ,   .          4                     state         <= waitingSvalid;5�_�   �   �           �   0   '    ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^�     �   /   1   6      *                     m_axis_tvalid <= '1';5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^�     �   .   0   7                              �   .   0   6    5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^0    �         7      0   type shiftState is (waitingSvalid, shifting);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^"�    �         8            �         7    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^"�     �         8      *      variable bitCounter :STD_LOGIC:='0';5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^"�    �         8      6      variable bitCounter :natural range 0 to 10:='0';5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%A     �               8   library IEEE;   use IEEE.STD_LOGIC_1164.ALL;       entity stretcher is       Port(     =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);   )           m_axis_tvalid : out STD_LOGIC;   )           m_axis_tlast  : out STD_LOGIC;   )           m_axis_tready : in  STD_LOGIC;       =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);   )           s_axis_tvalid : in  STD_LOGIC;   )           s_axis_tlast  : in  STD_LOGIC;   )           s_axis_tready : out STD_LOGIC;       )           clk           : in  STD_LOGIC;   *           rst           : in  STD_LOGIC);   end stretcher;       'architecture Behavioral of stretcher is   5   type shiftState is (waitingSvalid, waitingMready);   ,   signal state:shiftState := waitingSvalid;   begin          shift_reg:process (clk) is   7      variable bitCounter :natural range 0 to 10 :='0';      begin         if rising_edge(clk) then            if rst = '0' then   #            state <= waitingSvalid;            else               case state is   $               when waitingSvalid =>   '                  s_axis_tready <= '0';   -                  if s_axis_tvalid = '1' then   1                     state      <= waitingMready;   '                     bitCounter := '0';                     end if;   $               when waitingMready =>   -                  if m_axis_tready = '1' then   +                     if bitCounter < 8 then   /                        m_axis_tvalid   <= '1';   D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);   8                        bitCounter      := bitCounter+1;                        else   7                        state         <= waitingSvalid;   +                        s_axis_tready <= 1;                        end if;                     else   *                     m_axis_tvalid <= '0';                     end if;               end case;         end if;      end process shift_reg;       end Behavioral;5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%Z     �   4   6                end if;5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%z     �   5   7             end process shift_reg;5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%�     �   4   6   8    �   5   6   8    5�_�   �   �           �   6   	    ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%�     �   5   7                   end if;5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            .           /           V        ^%�    �   6   8                end process shift_reg;5�_�   �   �           �   /   )    ����                                                                                                                                                                                                                                                                                                                                                             ^2�     �   .   0   9      +                        s_axis_tready <= 1;5�_�   �   �   �       �   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^2�    �   .   0   9      ,                        s_axis_tready <= '1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^3M   	 �         9      7      variable bitCounter :natural range 0 to 10 :='0';5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                               0          5       v   5    ^3�   
 �         9      7      variable bitCounter :integer range 0 to 10 :='0';5�_�   �   �           �   %   #    ����                                                                                                                                                                                                                                                                                                                                                             ^3�     �   $   &   9      '                     bitCounter := '0';5�_�   �   �           �   %   $    ����                                                                                                                                                                                                                                                                                                                                                             ^3�    �   $   &   9      &                     bitCounter := 0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^8�     �          9    �          9    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^8�     �                 '                  s_axis_tready <= '0';5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^8�    �   7   9   :         end process shift_reg;�   6   8   :            end if;�   5   7   :               end if;�   4   6   :                  end case;�   3   5   :                        end if;�   2   4   :      *                     m_axis_tvalid <= '0';�   1   3   :                        else�   0   2   :                           end if;�   /   1   :      -                        s_axis_tready <= '1';�   .   0   :      7                        state         <= waitingSvalid;�   -   /   :                           else�   ,   .   :      8                        bitCounter      := bitCounter+1;�   +   -   :      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   :      /                        m_axis_tvalid   <= '1';�   )   +   :      +                     if bitCounter < 8 then�   (   *   :      -                  if m_axis_tready = '1' then�   '   )   :      $               when waitingMready =>�   &   (   :                        end if;�   %   '   :      %                     bitCounter := 0;�   $   &   :      1                     state      <= waitingMready;�   #   %   :      -                  if s_axis_tvalid = '1' then�   "   $   :      '                  s_axis_tready <= '0';�   !   #   :      $               when waitingSvalid =>�       "   :                  case state is�      !   :               else�          :      !            s_axis_tready <= '0';�         :      +            state         <= waitingSvalid;�         :               if rst = '0' then�         :            if rising_edge(clk) then�         :         begin�         :      1      variable bitCounter :integer range 0 to 10;�         :         shift_reg:process (clk) is�         :      ,   signal state:shiftState := waitingSvalid;�         :      5   type shiftState is (waitingSvalid, waitingMready);�         :      *           rst           : in  STD_LOGIC);�         :      )           clk           : in  STD_LOGIC;�         :      )           s_axis_tready : out STD_LOGIC;�         :      )           s_axis_tlast  : in  STD_LOGIC;�         :      )           s_axis_tvalid : in  STD_LOGIC;�   
      :      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   :      )           m_axis_tready : in  STD_LOGIC;�      	   :      )           m_axis_tlast  : out STD_LOGIC;�         :      )           m_axis_tvalid : out STD_LOGIC;�         :      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         :          Port(  �                #            state <= waitingSvalid;�                 !            s_axis_tready <= '0';5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                                                V       ^9r     �   /   1   :    �   0   1   :    5�_�   �   �           �   0   ,    ����                                                                                                                                                                                                                                                                                                                                                V       ^9t     �   /   1   ;      /                        m_axis_tvalid   <= '1';5�_�   �   �   �       �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9{     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      0                        s_axis_tready <= '   1';�   /   1   ;      0                        m_axis_tvalid   <= ' 0';�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   .   0          7                        state         <= waitingSvalid;�   0   2          -                        s_axis_tready <= '1';�   /   1          /                        m_axis_tvalid   <= '0';5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9~     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      0                        s_axis_tready <= '   1';�   /   1   ;      0                        m_axis_tvalid   <= ' 0';�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   .   0          7                        state         <= waitingSvalid;�   0   2          0                        s_axis_tready <= '   1';�   /   1          0                        m_axis_tvalid   <= ' 0';5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      7                        s_axis_tready <= '   1'       ;�   /   1   ;      7                        m_axis_tvalid   <= ' 0'       ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   0   2          0                        s_axis_tready <= '   1';�   /   1          0                        m_axis_tvalid   <= ' 0';�   .   0          7                        state         <= waitingSvalid;5�_�   �   �   �       �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      7                        s_axis_tready <= '   1'       ;�   /   1   ;      7                        m_axis_tvalid   <= ' 0'       ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   .   0          7                        state         <= waitingSvalid;�   0   2          7                        s_axis_tready <= '   1'       ;�   /   1          7                        m_axis_tvalid   <= ' 0'       ;5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      /                        s_axis_tready <= ' 1' ;�   /   1   ;      /                        m_axis_tvalid <= ' 0' ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   0   2          7                        s_axis_tready <= '   1'       ;�   /   1          7                        m_axis_tvalid   <= ' 0'       ;�   .   0          7                        state         <= waitingSvalid;5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      /                        s_axis_tready <= ' 1' ;�   /   1   ;      /                        m_axis_tvalid <= ' 0' ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   .   0          7                        state         <= waitingSvalid;�   0   2          /                        s_axis_tready <= ' 1' ;�   /   1          /                        m_axis_tvalid <= ' 0' ;5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      7                        s_axis_tready <= ' 1'         ;�   /   1   ;      7                        m_axis_tvalid <= ' 0'         ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   0   2          /                        s_axis_tready <= ' 1' ;�   /   1          /                        m_axis_tvalid <= ' 0' ;�   .   0          7                        state         <= waitingSvalid;5�_�   �   �           �   0   *    ����                                                                                                                                                                                                                                                                                                                            0   *       1   *          *    ^9�     �   /   2   ;      7                        m_axis_tvalid <= ' 0'         ;   7                        s_axis_tready <= ' 1'         ;5�_�   �   �   �       �   /        ����                                                                                                                                                                                                                                                                                                                            /   *       1   *       V   *    ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      7                        s_axis_tready <= ' 1'         ;�   /   1   ;      7                        m_axis_tvalid <= ' 0'         ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   .   0          7                        state         <= waitingSvalid;�   0   2          6                        s_axis_tready <= '1'         ;�   /   1          6                        m_axis_tvalid <= '0'         ;5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /   *       1   *       V   *    ^9�     �   8   :   ;         end process shift_reg;�   7   9   ;            end if;�   6   8   ;               end if;�   5   7   ;                  end case;�   4   6   ;                        end if;�   3   5   ;      *                     m_axis_tvalid <= '0';�   2   4   ;                        else�   1   3   ;                           end if;�   0   2   ;      /                        s_axis_tready <= ' 1' ;�   /   1   ;      /                        m_axis_tvalid <= ' 0' ;�   .   0   ;      7                        state         <= waitingSvalid;�   -   /   ;                           else�   ,   .   ;      8                        bitCounter      := bitCounter+1;�   +   -   ;      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   *   ,   ;      /                        m_axis_tvalid   <= '1';�   )   +   ;      +                     if bitCounter < 8 then�   (   *   ;      -                  if m_axis_tready = '1' then�   '   )   ;      $               when waitingMready =>�   &   (   ;                        end if;�   %   '   ;      %                     bitCounter := 0;�   $   &   ;      1                     state      <= waitingMready;�   #   %   ;      -                  if s_axis_tvalid = '1' then�   "   $   ;      '                  s_axis_tready <= '0';�   !   #   ;      $               when waitingSvalid =>�       "   ;                  case state is�      !   ;               else�          ;      !            s_axis_tready <= '0';�         ;      +            state         <= waitingSvalid;�         ;               if rst = '0' then�         ;            if rising_edge(clk) then�         ;         begin�         ;      1      variable bitCounter :integer range 0 to 10;�         ;         shift_reg:process (clk) is�         ;      ,   signal state:shiftState := waitingSvalid;�         ;      5   type shiftState is (waitingSvalid, waitingMready);�         ;      *           rst           : in  STD_LOGIC);�         ;      )           clk           : in  STD_LOGIC;�         ;      )           s_axis_tready : out STD_LOGIC;�         ;      )           s_axis_tlast  : in  STD_LOGIC;�         ;      )           s_axis_tvalid : in  STD_LOGIC;�   
      ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   ;      )           m_axis_tready : in  STD_LOGIC;�      	   ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�         ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         ;          Port(  �   0   2          7                        s_axis_tready <= ' 1'         ;�   /   1          7                        m_axis_tvalid <= ' 0'         ;�   .   0          7                        state         <= waitingSvalid;5�_�   �   �           �   0   *    ����                                                                                                                                                                                                                                                                                                                            0   *       1   *          *    ^9�     �   /   2   ;      /                        m_axis_tvalid <= ' 0' ;   /                        s_axis_tready <= ' 1' ;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            0   *       1   *          *    ^9�     �      !   ;    �       !   ;    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            1   *       2   *          *    ^9�     �      !          .                        m_axis_tvalid <= '0' ;5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                 V       ^9�     �   9   ;   <         end process shift_reg;�   8   :   <            end if;�   7   9   <               end if;�   6   8   <                  end case;�   5   7   <                        end if;�   4   6   <      *                     m_axis_tvalid <= '0';�   3   5   <                        else�   2   4   <                           end if;�   1   3   <      .                        s_axis_tready <= '1' ;�   0   2   <      .                        m_axis_tvalid <= '0' ;�   /   1   <      7                        state         <= waitingSvalid;�   .   0   <                           else�   -   /   <      8                        bitCounter      := bitCounter+1;�   ,   .   <      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   +   -   <      /                        m_axis_tvalid   <= '1';�   *   ,   <      +                     if bitCounter < 8 then�   )   +   <      -                  if m_axis_tready = '1' then�   (   *   <      $               when waitingMready =>�   '   )   <                        end if;�   &   (   <      %                     bitCounter := 0;�   %   '   <      1                     state      <= waitingMready;�   $   &   <      -                  if s_axis_tvalid = '1' then�   #   %   <      '                  s_axis_tready <= '0';�   "   $   <      $               when waitingSvalid =>�   !   #   <                  case state is�       "   <               else�      !   <      #            m_axis_tvalid <= ' 0' ;�          <      "            s_axis_tready <= ' 0';�         <      +            state         <= waitingSvalid;�         <               if rst = '0' then�         <            if rising_edge(clk) then�         <         begin�         <      1      variable bitCounter :integer range 0 to 10;�         <         shift_reg:process (clk) is�         <      ,   signal state:shiftState := waitingSvalid;�         <      5   type shiftState is (waitingSvalid, waitingMready);�         <      *           rst           : in  STD_LOGIC);�         <      )           clk           : in  STD_LOGIC;�         <      )           s_axis_tready : out STD_LOGIC;�         <      )           s_axis_tlast  : in  STD_LOGIC;�         <      )           s_axis_tvalid : in  STD_LOGIC;�   
      <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   <      )           m_axis_tready : in  STD_LOGIC;�      	   <      )           m_axis_tlast  : out STD_LOGIC;�         <      )           m_axis_tvalid : out STD_LOGIC;�         <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         <          Port(  �                +            state         <= waitingSvalid;�      !          "            m_axis_tvalid <= '0' ;�                 !            s_axis_tready <= '0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^9�     �      !   <      "            s_axis_tready <= ' 0';   #            m_axis_tvalid <= ' 0' ;5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                                                        ^9�    �      !   <      "            m_axis_tvalid <= '0' ;5�_�   �   �   �       �            ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;E     �       "   <    5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;F     �       "   =       �   !   "   =    5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;H     �       "          m_axis_tdata_tb5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;K     �       "   =                  m_axis_tdata_tb5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;L     �       #   =                  m_axis_tdata5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;Z     �       "   >      %            m_axis_tdata <= (others=>5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;b    �   !   "           5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                            !   
          
       V   
    ^;h    �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      *                     m_axis_tvalid <= '0';�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      .                        s_axis_tready <= '1' ;�   1   3   =      .                        m_axis_tvalid <= '0' ;�   0   2   =      7                        state         <= waitingSvalid;�   /   1   =                           else�   .   0   =      8                        bitCounter      := bitCounter+1;�   -   /   =      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   ,   .   =      /                        m_axis_tvalid   <= '1';�   +   -   =      +                     if bitCounter < 8 then�   *   ,   =      -                  if m_axis_tready = '1' then�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      %                     bitCounter := 0;�   &   (   =      1                     state      <= waitingMready;�   %   '   =      -                  if s_axis_tvalid = '1' then�   $   &   =      '                  s_axis_tready <= '0';�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      1      variable bitCounter :integer range 0 to 10;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �                +            state         <= waitingSvalid;�       "          *            m_axis_tdata <= (others=>'0');�      !          !            m_axis_tvalid <= '0';�                 !            s_axis_tready <= '0';5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            %   %       %   %       V   %    ^C�     �   $   %          '                  s_axis_tready <= '0';5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            %   %       %   %       V   %    ^C�     �   %   '   <    �   &   '   <    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            %   %       %   %       V   %    ^C�     �   %   '          '                  s_axis_tready <= '0';5�_�   �   �   �       �   &        ����                                                                                                                                                                                                                                                                                                                            &          (          V       ^C�     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      *                     m_axis_tvalid <= '0';�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      .                        s_axis_tready <= '1' ;�   1   3   =      .                        m_axis_tvalid <= '0' ;�   0   2   =      7                        state         <= waitingSvalid;�   /   1   =                           else�   .   0   =      8                        bitCounter      := bitCounter+1;�   -   /   =      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   ,   .   =      /                        m_axis_tvalid   <= '1';�   +   -   =      +                     if bitCounter < 8 then�   *   ,   =      -                  if m_axis_tready = '1' then�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      *                     bitCounter :=      0;�   &   (   =      1                     state      <= waitingMready;�   %   '   =      +                     s_axis_tready <= ' 0';�   $   &   =      -                  if s_axis_tvalid = '1' then�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      1      variable bitCounter :integer range 0 to 10;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   %   '          *                     s_axis_tready <= '0';�   '   )          %                     bitCounter := 0;5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            &           (           V        ^C�     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      *                     m_axis_tvalid <= '0';�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      .                        s_axis_tready <= '1' ;�   1   3   =      .                        m_axis_tvalid <= '0' ;�   0   2   =      7                        state         <= waitingSvalid;�   /   1   =                           else�   .   0   =      8                        bitCounter      := bitCounter+1;�   -   /   =      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   ,   .   =      /                        m_axis_tvalid   <= '1';�   +   -   =      +                     if bitCounter < 8 then�   *   ,   =      -                  if m_axis_tready = '1' then�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      *                     bitCounter :=      0;�   &   (   =      1                     state      <= waitingMready;�   %   '   =      +                     s_axis_tready <= ' 0';�   $   &   =      -                  if s_axis_tvalid = '1' then�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      1      variable bitCounter :integer range 0 to 10;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   %   '          +                     s_axis_tready <= ' 0';�   '   )          *                     bitCounter :=      0;5�_�   �   �   �       �   &        ����                                                                                                                                                                                                                                                                                                                            &           (           V        ^C�     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      *                     m_axis_tvalid <= '0';�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      .                        s_axis_tready <= '1' ;�   1   3   =      .                        m_axis_tvalid <= '0' ;�   0   2   =      7                        state         <= waitingSvalid;�   /   1   =                           else�   .   0   =      8                        bitCounter      := bitCounter+1;�   -   /   =      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);�   ,   .   =      /                        m_axis_tvalid   <= '1';�   +   -   =      +                     if bitCounter < 8 then�   *   ,   =      -                  if m_axis_tready = '1' then�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      (                     bitCounter    := 0;�   &   (   =      4                     state         <= waitingMready;�   %   '   =      +                     s_axis_tready <= ' 0';�   $   &   =      -                  if s_axis_tvalid = '1' then�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      1      variable bitCounter :integer range 0 to 10;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   %   '          +                     s_axis_tready <= ' 0';�   &   (          1                     state      <= waitingMready;�   '   )          *                     bitCounter :=      0;5�_�   �   �           �   &   '    ����                                                                                                                                                                                                                                                                                                                            &           (           V        ^C�     �   %   '   =      +                     s_axis_tready <= ' 0';5�_�   �   �           �      .    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^C�    �         =      1      variable bitCounter :integer range 0 to 10;5�_�   �   �           �   &   '    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^K     �   %   '   =      *                     s_axis_tready <= '0';5�_�   �              �   +   '    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^K     �   *   ,   =    �   +   ,   =    5�_�   �                +   '    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^K     �   *   ,   >      *                     s_axis_tready <= '1';5�_�                  4       ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^KK    �   3   4          .                        s_axis_tready <= '1' ;5�_�                 %   -    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M?     �   $   &   =      -                  if s_axis_tvalid = '1' then5�_�                 &   *    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^ML     �   %   '   =      *                     s_axis_tready <= '1';5�_�                 '   4    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^MT     �   &   (   =      4                     state         <= waitingMready;5�_�                 +   *    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^Ma     �   *   ,   =      *                     s_axis_tready <= '0';5�_�                 ,   -    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^Mq     �   +   -   =      -                  if m_axis_tready = '1' then5�_�                 ,   5    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^Mv     �   +   -   =      5                  if m_axis_tready = '1' then      --5�_�    	             -   +    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   ,   .   =      +                     if bitCounter < 8 then5�_�    
          	   .   /    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   -   /   =      /                        m_axis_tvalid   <= '1';5�_�  	            
   /   D    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   .   0   =      D                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);5�_�  
               0   8    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   /   1   =      8                        bitCounter      := bitCounter+1;5�_�                 2   7    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   1   3   =      7                        state         <= waitingSvalid;5�_�                 3   .    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   2   4   =      .                        m_axis_tvalid <= '0' ;5�_�                 6   *    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   5   7   =      *                     m_axis_tvalid <= '0';5�_�                 6   �    ����                                                                                                                                                                                                                                                                                                                               .          /       v   /    ^M�     �   5   7   =      �                     m_axis_tvalid <= '0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito_5�_�               %   3    ����                                                                                                                                                                                                                                                                                                                            %   3       &   3          3    ^N	     �   %   '   =      T                     s_axis_tready <= '1';         --entonces yo tambien estoy listo�   $   &   =      ]                  if s_axis_tvalid = '1' then      --espero a que este listo para enviar algo5�_�                 '   6    ����                                                                                                                                                                                                                                                                                                                            %   3       &   3          3    ^N     �   &   (   =      p                     state         <= waitingMready;  --cambio de estado, y le doy un clk para que ponga el dato5�_�                 +   3    ����                                                                                                                                                                                                                                                                                                                            +   3       .   3          3    ^N     �   +   /   =      \                  if m_axis_tready = '1' then      --lo puedo empezar a mandar al otro lado?   Q                     if bitCounter < 8 then        --perfecto, porque bit voy?      _                        m_axis_tvalid   <= '1';    --como puedo mandar, le avoso que tengo dato�   *   ,   =      h                     s_axis_tready <= '0';         --el dato esta en la mesa, ya no quiero mas por ahora5�_�                 0   9    ����                                                                                                                                                                                                                                                                                                                            +   3       .   3          3    ^N     �   /   1   =      E                        bitCounter      := bitCounter+1; --incremento5�_�                 +   :    ����                                                                                                                                                                                                                                                                                                                            .   ;       +   ;       V   ;    ^N*     �   *   ,   =      q                     s_axis_tready <= '0';                  --el dato esta en la mesa, ya no quiero mas por ahora5�_�                 +   :    ����                                                                                                                                                                                                                                                                                                                            .   ;       +   ;       V   ;    ^N*     �   *   ,   =      p                     s_axis_tready <= '0';                 --el dato esta en la mesa, ya no quiero mas por ahora5�_�                 +   :    ����                                                                                                                                                                                                                                                                                                                            +   :       .   :       V   :    ^NF     �   *   ,   =      o                     s_axis_tready <= '0';                --el dato esta en la mesa, ya no quiero mas por ahora5�_�                  +   ;    ����                                                                                                                                                                                                                                                                                                                            +   ;       .   ;          ;    ^NI     �   +   /   =      e                  if m_axis_tready = '1' then               --lo puedo empezar a mandar al otro lado?   Z                     if bitCounter < 8 then                 --perfecto, porque bit voy?      h                        m_axis_tvalid   <= '1';             --como puedo mandar, le avoso que tengo dato�   *   ,   =      q                     s_axis_tready <= '0';                  --el dato esta en la mesa, ya no quiero mas por ahora5�_�    !            +        ����                                                                                                                                                                                                                                                                                                                            +   ;       -   ;       V   ;    ^NO     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      �                     m_axis_tvalid <= '0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      Z                        m_axis_tvalid <= '0' ;  --y aviso que no tengo mas nada que mandar�   1   3   =      ^                        state         <= waitingSvalid;  --termine de mandar, vuelvo a esperar�   0   2   =                           else�   /   1   =      H                        bitCounter      := bitCounter+1;    --incremento�   .   0   =      U                        m_axis_tdata(0) <= s_axis_tdata(bitCounter); --pongo el dato �   -   /   =      r                        m_axis_tvalid   <= '1';                       --como puedo mandar, le avoso que tengo dato�   ,   .   =      d                     if bitCounter < 8 then                           --perfecto, porque bit voy?   �   +   -   =      o                  if m_axis_tready = '1' then                         --lo puedo empezar a mandar al otro lado?�   *   ,   =      {                     s_axis_tready <= '0';                            --el dato esta en la mesa, ya no quiero mas por ahora�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      (                     bitCounter    := 0;�   &   (   =      v                     state         <= waitingMready;        --cambio de estado, y le doy un clk para que ponga el dato�   %   '   =      ]                     s_axis_tready <= '1';                  --entonces yo tambien estoy listo�   $   &   =      f                  if s_axis_tvalid = '1' then               --espero a que este listo para enviar algo�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  5�_�     "          !   +        ����                                                                                                                                                                                                                                                                                                                            /   0       +   0       V   0    ^NS     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      �                     m_axis_tvalid <= '0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      Z                        m_axis_tvalid <= '0' ;  --y aviso que no tengo mas nada que mandar�   1   3   =      ^                        state         <= waitingSvalid;  --termine de mandar, vuelvo a esperar�   0   2   =                           else�   /   1   =      H                        bitCounter      := bitCounter+1;    --incremento�   .   0   =      U                        m_axis_tdata(0) <= s_axis_tdata(bitCounter); --pongo el dato �   -   /   =      r                        m_axis_tvalid   <= '1';                       --como puedo mandar, le avoso que tengo dato�   ,   .   =      d                     if bitCounter < 8 then                           --perfecto, porque bit voy?   �   +   -   =      o                  if m_axis_tready = '1' then                         --lo puedo empezar a mandar al otro lado?�   *   ,   =      {                     s_axis_tready <= '0';                            --el dato esta en la mesa, ya no quiero mas por ahora�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      (                     bitCounter    := 0;�   &   (   =      v                     state         <= waitingMready;        --cambio de estado, y le doy un clk para que ponga el dato�   %   '   =      ]                     s_axis_tready <= '1';                  --entonces yo tambien estoy listo�   $   &   =      f                  if s_axis_tvalid = '1' then               --espero a que este listo para enviar algo�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  5�_�  !  #          "   +   E    ����                                                                                                                                                                                                                                                                                                                            +   E       .   E          E    ^NW     �   *   /   =      {                     s_axis_tready <= '0';                            --el dato esta en la mesa, ya no quiero mas por ahora   o                  if m_axis_tready = '1' then                         --lo puedo empezar a mandar al otro lado?   d                     if bitCounter < 8 then                           --perfecto, porque bit voy?      r                        m_axis_tvalid   <= '1';                       --como puedo mandar, le avoso que tengo dato5�_�  "  &          #   +   E    ����                                                                                                                                                                                                                                                                                                                            +   E       /   E          E    ^N[     �   +   0   =      n                  if m_axis_tready = '1' then                        --lo puedo empezar a mandar al otro lado?   c                     if bitCounter < 8 then                          --perfecto, porque bit voy?      q                        m_axis_tvalid   <= '1';                      --como puedo mandar, le avoso que tengo dato   U                        m_axis_tdata(0) <= s_axis_tdata(bitCounter); --pongo el dato �   *   ,   =      z                     s_axis_tready <= '0';                           --el dato esta en la mesa, ya no quiero mas por ahora5�_�  #  '  $      &   %   E    ����                                                                                                                                                                                                                                                                                                                            %   E       %   E       v   E    ^Nc     �   $   &   =      f                  if s_axis_tvalid = '1' then               --espero a que este listo para enviar algo5�_�  &  (          '   %        ����                                                                                                                                                                                                                                                                                                                            %   E       .   E       V   E    ^Nf     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      �                     m_axis_tvalid <= '0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   4   6   =                        else�   3   5   =                           end if;�   2   4   =      Z                        m_axis_tvalid <= '0' ;  --y aviso que no tengo mas nada que mandar�   1   3   =      ^                        state         <= waitingSvalid;  --termine de mandar, vuelvo a esperar�   0   2   =                           else�   /   1   =      H                        bitCounter      := bitCounter+1;    --incremento�   .   0   =      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   -   /   =      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   ,   .   =      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   +   -   =      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   *   ,   =      }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   )   +   =      $               when waitingMready =>�   (   *   =                        end if;�   '   )   =      (                     bitCounter    := 0;�   &   (   =      v                     state         <= waitingMready;        --cambio de estado, y le doy un clk para que ponga el dato�   %   '   =      ]                     s_axis_tready <= '1';                  --entonces yo tambien estoy listo�   $   &   =      f                  if s_axis_tvalid = '1' then               --espero e que este listo para enviar algo�   #   %   =      $               when waitingSvalid =>�   "   $   =                  case state is�   !   #   =               else�       "   =      -            m_axis_tdata  <= (others => '0');�      !   =      !            m_axis_tvalid <= '0';�          =      !            s_axis_tready <= '0';�         =      +            state         <= waitingSvalid;�         =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�      
   =      )           m_axis_tready : in  STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�         =      )           m_axis_tvalid : out STD_LOGIC;�         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  5�_�  '  )          (   %   <    ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^Nj     �   %   (   =      ]                     s_axis_tready <= '1';                  --entonces yo tambien estoy listo   v                     state         <= waitingMready;        --cambio de estado, y le doy un clk para que ponga el dato�   $   &   =      f                  if s_axis_tvalid = '1' then               --espero e que este listo para enviar algo5�_�  (  *          )   0   <    ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^Nn     �   /   1   =      H                        bitCounter      := bitCounter+1;    --incremento5�_�  )  +          *   2   9    ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^Nq     �   1   3   =      ^                        state         <= waitingSvalid;  --termine de mandar, vuelvo a esperar5�_�  *  ,          +   3   0    ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^Ns     �   2   4   =      Z                        m_axis_tvalid <= '0' ;  --y aviso que no tengo mas nada que mandar5�_�  +  -          ,   6   -    ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^Nv     �   5   7   =      �                     m_axis_tvalid <= '0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)5�_�  ,  .          -          ����                                                                                                                                                                                                                                                                                                                            %   <       '   <          <    ^N|     �         >       �         =    5�_�  -  /          .           ����                                                                                                                                                                                                                                                                                                                            (   <       *   <          <    ^N�     �                 5�_�  .  0          /      
    ����                                                                                                                                                                                                                                                                                                                            '   <       )   <          <    ^N�     �         ?      I--tomo 1 bute y mando 8 bytes en donde en cada uno de salida vale el bit05�_�  /              0      
    ����                                                                                                                                                                                                                                                                                                                            '   <       )   <          <    ^N�    �         @       �         ?    5�_�  #  %      &  $   %   E    ����                                                                                                                                                                                                                                                                                                                            /   E       %   E       V   E    ^N^     �   $   0   =      feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   veeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   }eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Xeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  $              %   %        ����                                                                                                                                                                                                                                                                                                                            /   E       %   E       V   E    ^N^     �   $   0   =      feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   veeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   }eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Xeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�                +        ����                                                                                                                                                                                                                                                                                                                            +   ;       -   ;       V   ;    ^NL     �   *   .   =      {eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   oeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�                   +        ����                                                                                                                                                                                                                                                                                                                            +   ;       -   ;       V   ;    ^NL     �   *   .   =      {eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   oeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�               %        ����                                                                                                                                                                                                                                                                                                                            %           &           V        ^N     �   $   '   =      ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�               %        ����                                                                                                                                                                                                                                                                                                                            6           %           V        ^M�     �   $   7   =      ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   peeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   heeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   \eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   _eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ueeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   ^eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Zeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeee   �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�               %        ����                                                                                                                                                                                                                                                                                                                            6           %           V        ^M�     �   '   )          9                     bitCounter    :=                  0;�   $   &          n                  if s_axis_tvalid = '                 1' then      --espero a que este listo para enviar algo�   %   '          d                     s_axis_tready <= '                1';         --entonces yo tambien estoy listo�   +   -          m                  if m_axis_tready = '                 1' then      --lo puedo empezar a mandar al otro lado?�   ,   .          _                     if bitCounter <                   8then        --perfecto, porque bit voy?�   -   /          j                        m_axis_tvalid   <= '           1';    --como puedo mandar, le avoso que tengo dato�   .   0          f                        m_axis_tdata(                  0) <= s_axis_tdata(bitCounter); --pongo el dato�   /   1          F                        bitCounter      := bitCounter+ 1; --incremento�   *   ,          x                     s_axis_tready <= '                0';         --el dato esta en la mesa, ya no quiero mas por ahora�   2   4          g                        m_axis_tvalid <= '             0' ;  --y aviso que no tengo mas nada que mandar�   5   7          �                     m_axis_tvalid <= '                0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�         =          Port(  �         =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tready : in  STD_LOGIC;�   
      =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           clk           : in  STD_LOGIC;�         =      *           rst           : in  STD_LOGIC);�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      ,   signal state:shiftState := waitingSvalid;�         =         shift_reg:process (clk) is�         =      0      variable bitCounter :integer range 0 to 8;�         =         begin�         =            if rising_edge(clk) then�         =               if rst = '0' then�         =      +            state         <= waitingSvalid;�          =      !            s_axis_tready <= '0';�      !   =      !            m_axis_tvalid <= '0';�       "   =      -            m_axis_tdata  <= (others => '0');�   !   #   =               else�   "   $   =                  case state is�   #   %   =      $               when waitingSvalid =>�   $   &   =      n                  if s_axis_tvalid = '                 1' then      --espero a que este listo para enviar algo�   %   '   =      d                     s_axis_tready <= '                1';         --entonces yo tambien estoy listo�   &   (   =      p                     state         <= waitingMready;  --cambio de estado, y le doy un clk para que ponga el dato�   '   )   =      9                     bitCounter    :=                  0;�   (   *   =                        end if;�   )   +   =      $               when waitingMready =>�   *   ,   =      x                     s_axis_tready <= '                0';         --el dato esta en la mesa, ya no quiero mas por ahora�   +   -   =      m                  if m_axis_tready = '                 1' then      --lo puedo empezar a mandar al otro lado?�   ,   .   =      _                     if bitCounter <                   8then        --perfecto, porque bit voy?�   -   /   =      j                        m_axis_tvalid   <= '           1';    --como puedo mandar, le avoso que tengo dato�   .   0   =      f                        m_axis_tdata(                  0) <= s_axis_tdata(bitCounter); --pongo el dato�   /   1   =      F                        bitCounter      := bitCounter+ 1; --incremento�   0   2   =                           else�   1   3   =      ^                        state         <= waitingSvalid;  --termine de mandar, vuelvo a esperar�   2   4   =      g                        m_axis_tvalid <= '             0' ;  --y aviso que no tengo mas nada que mandar�   3   5   =                           end if;�   4   6   =                        else�   5   7   =      �                     m_axis_tvalid <= '                0';   --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   6   8   =                        end if;�   7   9   =                  end case;�   8   :   =               end if;�   9   ;   =            end if;�   :   <   =         end process shift_reg;5�_�               %        ����                                                                                                                                                                                                                                                                                                                            6           %           V        ^M�     �   $   7   =      ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   peeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   heeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   \eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   _eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ueeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   ^eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Zeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeee   �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�               %        ����                                                                                                                                                                                                                                                                                                                            6           %           V        ^M�     �   $   7   =      ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   peeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   heeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   \eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   _eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ueeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   ^eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Zeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeee   �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�                 %        ����                                                                                                                                                                                                                                                                                                                            6           %           V        ^M�     �   $   7   =      ]eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   peeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   heeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   \eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   _eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ueeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeee   ^eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Zeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeee   �eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   &        ����                                                                                                                                                                                                                                                                                                                            &           (           V        ^C�     �   %   )   =      +eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   1eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �       �   �   �   &        ����                                                                                                                                                                                                                                                                                                                            &          (          V       ^C�     �   %   )   =      *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   1eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   %eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   &        ����                                                                                                                                                                                                                                                                                                                            &          (          V       ^C�     �   %   )   =      *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   1eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   %eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �      
    ����                                                                                                                                                                                                                                                                                                                            !   
          
       V   
    ^;e     �      "   =      +eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   !eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   !eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �            ����                                                                                                                                                                                                                                                                                                                                           	       V   	    ^;C     �       !   <    �      !   <      0 m_axis_tdata_tb           m_axis_tvalid <= '0';5�_�   �       �   �   �           ����                                                                                                                                                                                                                                                                                                                                                   V        ^9�     �      !   <      +eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   !eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   "eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �           ����                                                                                                                                                                                                                                                                                                                                                 V       ^9�     �      !   <      +eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   !eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   "eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   /        ����                                                                                                                                                                                                                                                                                                                            /   *       1   *       V   *    ^9�     �   .   2   ;      7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   6eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   6eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �       �   �   �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   .   2   ;      7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9�     �   .   2   ;      7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �       �   �   �   /        ����                                                                                                                                                                                                                                                                                                                            /           1           V        ^9y     �   .   2   ;      7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   /eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   -eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   /        ����                                                                                                                                                                                                                                                                                                                            /   ,       1   ,       V   ,    ^9v     �   .   2   ;      7eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   /eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   -eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   /   +    ����                                                                                                                                                                                                                                                                                                                                                             ^2�     �   .   0   9      -                        s_axis_tready <= '1';5�_�   �       �   �   �   )   &    ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^a     �   (   *   4      '                        m_axis_tvalid j5�_�   �           �   �   )        ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^]     �   (   +   4      -eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �      &    ����                                                                                                                                                                                                                                                                                                                                                  v       ^�     �         2      ,   signal state:shiftState := waitingSValid;5�_�   �           �   �   "       ����                                                                                                                                                                                                                                                                                                                                         "       v        ^�     �   !   #   2                         if  = '1' then5�_�   }              ~          ����                                                                                                                                                                                                                                                                                                                                         *       v   *    ^s     �         2    �         2      ,   signal state:shiftState := waitingS_Vali;5�_�   5           7   6           ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �          )    �          )       tateMealy_re        else5�_�                          ����                                                                                                                                                                                                                                                                                                                                                  V        ^v     �              5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         "         �         #         ooi5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^
�     �             �               !      if rising_byeedge(clk) then5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ^
m     �               >eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee       >eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   "eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee       #eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5��