Vim�UnDo� �զ&�c�~L��`�
��2/4A�?81�yy�   =                                   ^�    _�                              ����                                                                                                                                                                                                                                                                                                                                                             ^�    �                'architecture Behavioral of join_8to1 is�                end join_8to1;�                entity join_8to1 is5��