Vim�UnDo� �q��wq�����2���]�Mx�ZC�3���   ;   library IEEE;                          ^��   = _�                     &        ����                                                                                                                                                                                                                                                                                                                                                             ^�(     �   %   '   )    5�_�                    &        ����                                                                                                                                                                                                                                                                                                                                                             ^�)     �   &   (   *    �   &   '   *    5�_�                    &        ����                                                                                                                                                                                                                                                                                                                                                             ^�+     �   %   &           5�_�                    &       ����                                                                                                                                                                                                                                                                                                                                                             ^�/     �   %   '          ,                       misoSignal <= inData;5�_�                    &       ����                                                                                                                                                                                                                                                                                                                                                             ^�c     �   %   &          (                   misoSignal <= inData;5�_�                            ����                                                                                                                                                                                                                                                                                                                                      (          V       ^�r     �      )   )    �         )    5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^�y     �   (   *   >          process (clk)5�_�      	              )       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^�}     �   (   *   >          cs:process (clk)5�_�      
           	   )       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   (   *   >          cs:process (csj)5�_�   	              
   ,       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   +   -   >      $            if rising_edge(clk) then5�_�   
                 ,       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   +   -   >      %            if falling_edge(clk) then5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   +   -   >      $            if falling_edge(ck) then5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   )   *          0       variable count: integer range 0 to 8 :=0;5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            )          <          V       ^��     �   ,   .   =    �   -   .   =    5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   ,   .   >      ,                       misoSignal <= inData;5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   ,   .   >      +                      misoSignal <= inData;5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   ,   .   >      *                     misoSignal <= inData;5�_�                    +       ����                                                                                                                                                                                                                                                                                                                            )          =          V       ^��     �   *   ,   >      $            if falling_edge(cs) then5�_�                    .        ����                                                                                                                                                                                                                                                                                                                            .          2          V       ^��     �   -   .          D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;   0                    spi_miso   <= misoSignal(7);   +                    count      := count +1;   '                    if (count < 8) then   B                       misoSignal <= misoSignal(6 downto 0) & '0';5�_�                    .        ����                                                                                                                                                                                                                                                                                                                            .          2          V       ^��     �   -   .                              else   ,                       misoSignal <= inData;   G                       outData    <= mosiSignal(6 downto 0) & spi_mosi;   G                       ledsData   <= mosiSignal(2 downto 0) & spi_mosi;   '                       count      := 0;5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^��     �   -   /                              end if;5�_�                    /        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   .   /                          else                       count := 0;                   end if;5�_�                    /       ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^��     �   .   0                       end if;5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^��    �         1          process (clk)5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^��     �   (   *   1          cs:process (cs)5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^��     �         1          spi:process (clk)5�_�                           ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^��    �         1          spi_prox:process (clk)5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            )          0                 ^�    �   )   1   1              begin   #            if rising_edge(cs) then   "                if (cs = '0') then   )                    misoSignal <= inData;                    end if;                 end if;           end process;�   (   *   1          cs_proc:process (cs)5�_�                    )       ����                                                                                                                                                                                                                                                                                                                            )          0                 ^�(     �   (   1   1       --   cs_proc:process (cs)    --       begin   % --           if rising_edge(cs) then   $ --               if (cs = '0') then   + --                   misoSignal <= inData;    --                end if;    --             end if;    --       end process;5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                            )          0                 ^��     �   +   ,          "                if (cs = '0') then5�_�                     -       ����                                                                                                                                                                                                                                                                                                                            )          /                 ^��     �   ,   -                           end if;5�_�      !               -       ����                                                                                                                                                                                                                                                                                                                            )          .                 ^��     �   ,   .                        end if;5�_�       "           !   -       ����                                                                                                                                                                                                                                                                                                                            )          .                 ^��     �   ,   .   /                       end if;5�_�   !   #           "   -       ����                                                                                                                                                                                                                                                                                                                            )          .                 ^��     �   ,   .   /                    end if;5�_�   "   $           #   +       ����                                                                                                                                                                                                                                                                                                                            )          .                 ^��    �   *   ,          #            if rising_edge(cs) then5�_�   #   %           $   ,       ����                                                                                                                                                                                                                                                                                                                            )          .                 ^��    �   +   -          )                    misoSignal <= inData;5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             ^�'     �         /          spi_proc:process (clk)5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             ^�9     �         /    �         /    5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             ^�<     �         0      $            if rising_edge(clk) then5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             ^�F     �         0    �         0    5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             ^�I     �                ,                       misoSignal <= inData;5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             ^�J     �         2                     �         1    5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             ^�d     �         2      #            if rising_edge(cs) then5�_�   +   /           ,   ,        ����                                                                                                                                                                                                                                                                                                                            ,           1                   ^��    �   ,   2   2              begin   "           if rising_edge(cs) then   #              misoSignal <= inData;              end if;           end process;�   +   -   2          cs_proc:process (cs)5�_�   ,   0   -       /   *       ����                                                                                                                                                                                                                                                                                                                            ,           1                   ^��     �   )   +   2    �   *   +   2    5�_�   /   1           0   +       ����                                                                                                                                                                                                                                                                                                                            -           2                   ^��    �   *   ,                       end if;5�_�   0   2           1   -        ����                                                                                                                                                                                                                                                                                                                            -           2           V        ^   
 �   ,   -          --    cs_proc:process (cs)   --        begin   $--           if rising_edge(cs) then   %--              misoSignal <= inData;   --           end if;   --        end process;5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^��    �         -          spi_proc:process (clk,cs)5�_�   2   4           3   '       ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^�    �   &   (                          else 5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^�E     �         -                  else5�_�   4   6           5   +   
    ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^�S    �   *   +                    end if;5�_�   5   7           6   $   %    ����                                                                                                                                                                                                                                                                                                                                                             ^�(     �   #   %   ,      G                       ledsData   <= mosiSignal(2 downto 0) & spi_mosi;5�_�   6   8           7   $   5    ����                                                                                                                                                                                                                                                                                                                                                             ^�/    �   #   %   ,      L                       ledsData   <= cs & mosiSignal(2 downto 0) & spi_mosi;5�_�   7   9           8   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^�w     �   +   -   ,    �   ,            5�_�   8   :           9   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^�x     �   +   -          L                       ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   9   ;           :   $       ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   #   %   -      L                       ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   :   <           ;   ,   &    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   +   -   -      =        ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   ;   =           <   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   +   -   -      =        ledsData   <= cs & mosiSignal(2 downto 0) & spi_mosi;5�_�   <   >           =   ,   .    ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   +   -   -      :        ledsData   <= cs & outData(2 downto 0) & spi_mosi;5�_�   =   ?           >   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   +   -   -      /        ledsData   <= cs & outData(2 downto 0);5�_�   >   @           ?   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   +   -   -      3        ledsData   <= not cs & outData(2 downto 0);5�_�   ?   A           @   ,        ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �               -   library IEEE;   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.NUMERIC_STD.ALL;       entity spi28b is   &    Port ( spi_mosi : in    STD_LOGIC;   &           spi_miso : out   STD_LOGIC;   &           cs       : in    std_logic;   :           outData  : out   std_logic_vector (7 downto 0);   :           inData   : in    std_logic_vector (7 downto 0);   :           ledsData : out   std_logic_vector (3 downto 0);   '           clk      : in    STD_LOGIC);   end spi28b;       $architecture Behavioral of spi28b is   I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');   I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');       begin         spi_proc:process (clk,cs) is   0       variable count: integer range 0 to 8 :=0;           begin   $            if falling_edge(cs) then   $               misoSignal <= inData;               end if;   $            if rising_edge(clk) then   "                if (cs = '0') then   D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;   0                    spi_miso   <= misoSignal(7);   +                    count      := count +1;   '                    if (count < 8) then   B                       misoSignal <= misoSignal(6 downto 0) & '0';                       else   ,                       misoSignal <= inData;   G                       outData    <= mosiSignal(6 downto 0) & spi_mosi;   N                       --ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;   '                       count      := 0;                       end if;                    else                       count := 0;                   end if;                end if;           end process;   6        ledsData   <= not cs & mosiSignal(2 downto 0);   end Behavioral;5�_�   @   B           A   $       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      N                       --ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   A   C           B   $       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      M                       -ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   B   D           C   $       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      L                       ledsData   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   C   E           D   $   1    ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      X                       ledsData(2 downto 0)   <= cs & mosiSignal(1 downto 0) & spi_mosi;5�_�   D   F           E   $   1    ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      W                       ledsData(2 downto 0)   <= s & mosiSignal(1 downto 0) & spi_mosi;5�_�   E   G           F   $   1    ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      V                       ledsData(2 downto 0)   <=  & mosiSignal(1 downto 0) & spi_mosi;5�_�   F   H           G   $   1    ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      U                       ledsData(2 downto 0)   <= & mosiSignal(1 downto 0) & spi_mosi;5�_�   G   I           H   $   1    ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   #   %   .      T                       ledsData(2 downto 0)   <=  mosiSignal(1 downto 0) & spi_mosi;5�_�   H   J           I   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   +   -   .               ledsData(3)   <= not cs;5�_�   I   K           J   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   +   -   .              ledsData(3)   <= ot cs;5�_�   J   L           K   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   +   -   .              ledsData(3)   <= t cs;5�_�   K   M           L   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   +   -   .              ledsData(3)   <=  cs;5�_�   L   N           M   -       ����                                                                                                                                                                                                                                                                                                                                                             ^	��    �   ,   -          7        ledsData(2 downto 0) <= mosiSignal(2 downto 0);5�_�   M   O           N   "        ����                                                                                                                                                                                                                                                                                                                                                             ^	ϥ    �   !   #   -      ,                       misoSignal <= inData;5�_�   N   P           O   *       ����                                                                                                                                                                                                                                                                                                                                                             ^	�     �   )   +   .                      �   )   +   -    5�_�   O   Q           P           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �                $            if falling_edge(cs) then   $               misoSignal <= inData;               end if;5�_�   P   R           Q   '        ����                                                                                                                                                                                                                                                                                                                            '          '          V       ^	�!     �   &   *   *    �   '   (   *    �   &   '                       else if*5�_�   Q   S           R   '       ����                                                                                                                                                                                                                                                                                                                            '           )          V       ^	�#     �   &   )   -      $            if falling_edge(cs) then5�_�   R   T           S   )       ����                                                                                                                                                                                                                                                                                                                            '           *          V       ^	�&     �   (   *          $               misoSignal <= inData;5�_�   S   U           T   *       ����                                                                                                                                                                                                                                                                                                                            '           *          V       ^	�-     �   )   +   .    �   *   +   .    5�_�   T   V           U   *       ����                                                                                                                                                                                                                                                                                                                            '           +          V       ^	�.    �   )   +                      end if;5�_�   U   W           V   +       ����                                                                                                                                                                                                                                                                                                                            '           +          V       ^	�9    �   *   +                      end if;5�_�   V   X           W   +       ����                                                                                                                                                                                                                                                                                                                            '           +          V       ^	�;     �   *   ,                       end if;5�_�   W   Y           X   '        ����                                                                                                                                                                                                                                                                                                                            '          +          V       ^	�J     �   &   ,   .                      else   +                   if falling_edge(cs) then   +                      misoSignal <= inData;                      end if;                   end if;5�_�   X   Z           Y   '       ����                                                                                                                                                                                                                                                                                                                            '          +                 ^	�Q     �   &   ,   .                   else   (                if falling_edge(cs) then   (                   misoSignal <= inData;                   end if;                end if;5�_�   Y   [           Z   '       ����                                                                                                                                                                                                                                                                                                                            '          +                 ^	�R     �   &   (                      else5�_�   Z   `           [   (        ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	�V    �   *   ,                      end if;�   )   +                         end if;�   (   *          '                  misoSignal <= inData;�   '   )          '               if falling_edge(cs) then5�_�   [   a   ^       `          ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	�4    �         .      0       variable count: integer range 0 to 8 :=0;5�_�   `   b           a      -    ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	�h     �         .      0                    spi_miso   <= misoSignal(7);5�_�   a   c           b      2    ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	�i     �         .      5                    spi_miso   <= misoSignal(count7);5�_�   b   d           c           ����                                                                                                                                                                                                                                                                                                                               2          2       V   2    ^	�j     �                4                    spi_miso   <= misoSignal(count);5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                               2          2       V   2    ^	�l    �         -    �         -    5�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�o     �                +                    count      := count +1;5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�o    �         -    �         -    5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�x     �                +                    count      := count +1;5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�z    �         -    �         -    5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                                                V       ^	ؘ    �         .      B                       misoSignal <= misoSignal(6 downto 0) & '0';5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                                                V       ^	؟     �         .      '                    if (count < 8) then5�_�   j   l           k           ����                                                                                                                                                                                                                                                                                                                                                V       ^	أ   ! �         .                          else5�_�   k   m           l           ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �                D                    --   misoSignal <= misoSignal(6 downto 0) & '0';   --                    else   .--                       misoSignal <= inData;5�_�   l   n           m   $       ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �   #   $                       else5�_�   m   o           n   $        ����                                                                                                                                                                                                                                                                                                                            $          &          V       ^	��     �   #   $          (                if falling_edge(cs) then   (                   misoSignal <= inData;                   end if;5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ^	��     �         '    �         '    5�_�   o   q           p           ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �         *    �         *    5�_�   p   r           q          ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �         -         spi_proc:process (clk,cs) is5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -         cs_proc:process (clk,cs) is5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -         cs_proc:process (lk,cs) is5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -         cs_proc:process (k,cs) is5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -         cs_proc:process (,cs) is5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �                0       variable count: natural range 0 to 8 :=0;5�_�   v   x           w           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�	     �                                end if;�                (                   misoSignal <= inData;�                (                if falling_edge(cs) then5�_�   w   y           x          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         ,    �         ,    5�_�   x   z           y          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �                0       variable count: natural range 0 to 8 :=0;5�_�   y   {           z          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -                 �         ,    5�_�   z   |           {          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         -    5�_�   {   }           |          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�      �         .         spi_proc:process (clk,cs) is5�_�   |   ~           }          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�      �         .         spi_proc:process (clkcs) is5�_�   }              ~          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�      �         .         spi_proc:process (clks) is5�_�   ~   �              $        ����                                                                                                                                                                                                                                                                                                                            $          &          V       ^	�;   " �   ,   .   .              ledsData(3)   <= cs;�   +   -   .              end process;�   *   ,   .                   end if;�   )   +   .                      end if;�   (   *   .                         count := 0;�   '   )   .                       else �   &   (   .                          end if;�   %   '   .      1                       count                := 0;�   $   &   .      Q                       ledsData(2 downto 0) <= mosiSignal(1 downto 0) & spi_mosi;�   #   %   .      Q                       outData              <= mosiSignal(6 downto 0) & spi_mosi;�   "   $   .      '                    if (count = 8) then�   !   #   .      +                    count      := count +1;�       "   .      4                    spi_miso   <= misoSignal(count);�      !   .      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�          .      "                if (cs = '0') then�         .      $            if rising_edge(clk) then�         .              begin�         .      0       variable count: natural range 0 to 8 :=0;�         .         spi_proc:process (clk) is�         .              end process cs_proc;�         .                 end if;�         .      #              misoSignal <= inData;�         .      #           if falling_edge(cs) then�         .              begin�         .         cs_proc:process (cs) is�         .      begin   �         .      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         .      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         .      '           clk      : in    STD_LOGIC);�   
      .      :           ledsData : out   std_logic_vector (3 downto 0);�   	      .      :           inData   : in    std_logic_vector (7 downto 0);�      
   .      :           outData  : out   std_logic_vector (7 downto 0);�      	   .      &           cs       : in    std_logic;�         .      &           spi_miso : out   STD_LOGIC;�         .      &    Port ( spi_mosi : in    STD_LOGIC;�   #   %          G                       outData    <= mosiSignal(6 downto 0) & spi_mosi;�   %   '          '                       count      := 0;�   $   &          S                       ledsData(2 downto 0)   <= mosiSignal(1 downto 0) & spi_mosi;5�_�      �           �   !   -    ����                                                                                                                                                                                                                                                                                                                            $          &          V       ^	�&   # �       "   .      4                    spi_miso   <= misoSignal(count);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $          &          V       ^	��     �         .      0       variable count: natural range 0 to 8 :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $          &          V       ^	��     �         .         spi_proc:process (clk) is5�_�   �   �           �   ,        ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �   +   /   .    �   ,   -   .    5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �   ,   .   1    �   -   .   1    5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                                                V       ^	��     �   ,   .   2                         count := 0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                          ^	��     �         2              begin   #           if falling_edge(cs) then   #              misoSignal <= inData;              end if;           end process cs_proc;�         2         cs_proc:process (cs) is5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                        ^	��   $ �         2      //   cs_proc:process (cs) is   //        begin   %//           if falling_edge(cs) then   %//              misoSignal <= inData;   //           end if;   //        end process cs_proc;5�_�   �   �           �   -        ����                                                                                                                                                                                                                                                                                                                            .   "       -          V   "    ^	�u   % �   0   2   2              ledsData(3)   <= cs;�   /   1   2              end process;�   .   0   2                 end if;�   -   /   2      #              misoSignal <= inData;�   ,   .   2                    count      := 0;�   +   -   2      #           if falling_edge(cs) then�   *   ,   2                   end if;�   )   +   2                      end if;�   (   *   2                         count := 0;�   '   )   2                       else �   &   (   2                          end if;�   %   '   2      1                       count                := 0;�   $   &   2      Q                       ledsData(2 downto 0) <= mosiSignal(1 downto 0) & spi_mosi;�   #   %   2      Q                       outData              <= mosiSignal(6 downto 0) & spi_mosi;�   "   $   2      '                    if (count = 8) then�   !   #   2      +                    count      := count +1;�       "   2      6                    spi_miso   <= misoSignal(7-count);�      !   2      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�          2      "                if (cs = '0') then�         2      $            if rising_edge(clk) then�         2              begin�         2      0       variable count: integer range 0 to 8 :=0;�         2         spi_proc:process (clk,cs) is�         2      --        end process cs_proc;�         2      --           end if;�         2      %--              misoSignal <= inData;�         2      %--           if falling_edge(cs) then�         2      --        begin�         2      --   cs_proc:process (cs) is�         2      begin   �         2      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         2      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         2      '           clk      : in    STD_LOGIC);�   
      2      :           ledsData : out   std_logic_vector (3 downto 0);�   	      2      :           inData   : in    std_logic_vector (7 downto 0);�      
   2      :           outData  : out   std_logic_vector (7 downto 0);�      	   2      &           cs       : in    std_logic;�         2      &           spi_miso : out   STD_LOGIC;�         2      &    Port ( spi_mosi : in    STD_LOGIC;�   ,   .                        count := 0;�   -   /          #              misoSignal <= inData;5�_�   �   �   �       �   0        ����                                                                                                                                                                                                                                                                                                                            ,           /           V        ^	��     �   /   4   2    �   0   1   2    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            ,           /           V        ^	��     �   /   1   6      #           if falling_edge(cs) then5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            ,           /           V        ^	��     �   1   2          #              misoSignal <= inData;5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            0          0          v       ^	�     �   /   1   5      "           if rising_edge(cs) then5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            0          0          v       ^	�     �   /   1   5                 if cs) then5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            0          0          v       ^	�     �   /   1   5                 if cs = '1') then5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            0          0          v       ^	�     �   0   2   5                    count      := 0;5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^	�     �   '   (                           else                       count := 0;5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^	�   + �   *   +                        count      := 0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ^@�     �         2    �         2    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^@�     �         3      &           spi_miso : out   STD_LOGIC;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^@�     �         3      /           stop_dataspi_miso : out   STD_LOGIC;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      --   cs_proc:process (cs) is   --        begin   %--           if falling_edge(cs) then   %--              misoSignal <= inData;   --           end if;   --        end process cs_proc;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3         cs_proc:process (cs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3         s_proc:process (cs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3         _proc:process (cs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      '           clk      : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      +           spi_clk      : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      *           spi_clk     : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      )           spi_clk    : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      (           spi_clk   : in    STD_LOGIC);5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         3         spi_proc:process (clk,cs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �          3      $            if rising_edge(clk) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         3    �         3    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         4      '           spi_clk  : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         4      (           sspi_clk  : in    STD_LOGIC);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         4         stop_proc:process (cs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A$     �         5            �         4    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^A?     �         5      #           if falling_edge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AF     �         5      '           if rising_edge_edge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AF     �         5      &           if rising_edgeedge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AF     �         5      %           if rising_edgedge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AF     �         5      $           if rising_edgege(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AG     �         5      #           if rising_edgee(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AG     �         5      "           if rising_edge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AM     �         5      #              misoSignal <= inData;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AS     �                #              misoSignal <= inData;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^AT     �         6                    �         5    5�_�   �   �           �      #    ����                                                                                                                                                                                                                                                                                                                                                        ^A_     �         6      #              if counter = 100000005�_�   �   �           �      +    ����                                                                                                                                                                                                                                                                                                                                                        ^A�     �         9                       �         8    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                         ^A�     �      !   9              end process cs_proc;5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                         ^A�     �      !   9              end process ss_proc;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                         ^A�     �      !   9              end process s_proc;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                         ^A�   , �      !   9              end process _proc;5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                                                             ^A�   - �         9      '           spi_clk  : in    STD_LOGIC);5�_�   �   �           �      5    ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �         9      :      variable counter : integer range (0 to 10000000) :=05�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             ^A�   . �         9      9      variable counter : integer range (0 to 10000000 :=05�_�   �   �           �      8    ����                                                                                                                                                                                                                                                                                                                                                             ^A�   0 �         9      8      variable counter : integer range 0 to 10000000 :=05�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                             ^G6     �         9    �         9    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^G8     �         :      9      variable counter : integer range 0 to 10000000 :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^G<     �         :      8      signal  counter : integer range 0 to 10000000 :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^G@     �         :      ;      signal  stop_state : integer range 0 to 10000000 :=0;5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                               %          8       v   8    ^GE     �         :      =      signal  stop_state : STD_LOGIC range 0 to 10000000 :=0;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                               %          8       v   8    ^GL   1 �         :      ,                 stop_data <= not stop_data;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               %          8       v   8    ^GT     �         :      )      signal  stop_state : STD_LOGIC :=0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^GY     �                (      signal stop_state : STD_LOGIC :=0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^GZ     �         9    �         9    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^G[     �         :      (      signal stop_state : STD_LOGIC :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^G\   3 �         :      '     signal stop_state : STD_LOGIC :=0;5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                                                V       ^G�     �         :      &    signal stop_state : STD_LOGIC :=0;5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                V       ^G�   4 �         :      '    signal stop_state : STD_LOGIC :='0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^U
     �         :      -                 stop_data <= not stop_state;5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   :    �   "   #   :    5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      .                 stop_state <= not stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      %        stop_state <= not stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      $        stop_date <= not stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      #        stop_date <= ot stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      "        stop_date <= t stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;      !        stop_date <=  stop_state;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^U     �   !   #   ;               stop_date <= stop_state;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ^U"     �         ;      (              if counter = 10000000 then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ^U"     �         ;      '              if counter = 1000000 then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ^U#     �         ;      &              if counter = 100000 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^U$   5 �         ;      %              if counter = 10000 then5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                                                             ^V     �   9   ;   ;              ledsData(3)   <= cs;5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                                                             ^V!     �   -   /   ;      Q                       ledsData(2 downto 0) <= mosiSignal(1 downto 0) & spi_mosi;5�_�   �   �           �   .   :    ����                                                                                                                                                                                                                                                                                                                                                             ^V(   6 �   -   /   ;      Q                       ledsData(1 downto 0) <= mosiSignal(1 downto 0) & spi_mosi;5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                                                             ^W@     �   9   ;   ;      )        ledsData(3)   <= cs & stop_state;5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                                                             ^WB   7 �   9   ;   ;      )        ledsData(3)   <= cs ^ stop_state;5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                                                             ^WH   8 �   9   ;   ;      )        ledsData(3)   <= cs & stop_state;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^X     �         ;      $              if counter = 1000 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^X$     �         ;      (              if counter = 10000000 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^X'     �         ;      (              if counter = 60000000 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^X)   9 �         ;      (              if counter = 60000000 then5�_�   �              �      ,    ����                                                                                                                                                                                                                                                                                                                                                             ^Z*     �         ;      9      variable counter : integer range 0 to 10000000 :=0;5�_�   �                   ,    ����                                                                                                                                                                                                                                                                                                                                                             ^Z,   : �         ;      9      variable counter : integer range 0 to 60000000 :=0;5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             ^��     �         ;    �         ;    5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      &           stop_data: out   STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      -           start_rx_op_data: out   STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      ,           start_rx_p_data: out   STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      +           start_rx__data: out   STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      *           start_rx_data: out   STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      	   <      1           tx_laststart_rx_data: out   STD_LOGIC;5�_�    	                    ����                                                                                                                                                                                                                                                                                                                                         $       v   $    ^��     �      	   <      8           tx_paquet_laststart_rx_data: out   STD_LOGIC;5�_�    
          	          ����                                                                                                                                                                                                                                                                                                                                         $       v   $    ^��     �      	   <      ,           tx_paquet_lasta: out   STD_LOGIC;5�_�  	            
          ����                                                                                                                                                                                                                                                                                                                                         $       v   $    ^t   ; �                +           tx_paquet_last: out   STD_LOGIC;5�_�  
                       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �          ;      library IEEE;5�_�                         ����                                                                                                                                                                                                                                                                                                                                                             ^�   < �          ;      ribrary IEEE;5�_�                         ����                                                                                                                                                                                                                                                                                                                                                             ^��     �          ;      igibrary IEEE;5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             ^��   = �          ;      liibrary IEEE;5�_�   �           �   �           ����                                                                                                                                                                                                                                                                                                                                                         ^A�     �      !   9              end process ;5�_�   �       �   �   �          ����                                                                                                                                                                                                                                                                                                                                                        ^A     �         3      &           spi_clk : in    STD_LOGIC);5�_�   �   �       �   �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      &           spi_clk : in    STD_LOGIC);5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                                                        ^@�     �         3      %           spi_clk  in    STD_LOGIC);5�_�   �   �       �   �   -        ����                                                                                                                                                                                                                                                                                                                                                             ^	��   ' �   ,   .   2       --              count      := 0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                        ^	�     �         2         cs_proc:process (cs) is           begin   #           if falling_edge(cs) then   #              misoSignal <= inData;              end if;           end process cs_proc;5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                        ^	�     �         2                    �         3                    rst_count <= '1';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                        ^	��     �          3                     �      !   4      (               if (rst_count = '1') then   "                  rst_count = '0';                  end if5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                                        ^	��     �       "   6      #                  rst_count <= '0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         6                    rst_count <= '0';5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         6    �         6      #           if falling_edge(cs) then   #              misoSignal <= inData;                 rst_count <= '0';              end if;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         :      '           if rising_edge_edge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         :      "           if rising_edge(cs) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�     �         9                    rst_count <= '1';5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^	�"     �              5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                V       ^	�>     �   !   "   6                        �   !   #   7                        count := 0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�_     �         7         spi_proc:process (clkcs) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ^	�_     �         7         spi_proc:process (clks) is5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            -          .          V       ^	�_     �         7         spi_proc:process (clk) is5�_�   �   �           �   -        ����                                                                                                                                                                                                                                                                                                                            /          2          V       ^	�j     �   ,   /        5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^	�q     �   .   3        5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^	�w     �         1    �         1      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            0          0          V       ^	�y     �         2      H    signal rst_count : std_logic_vector (7 downto 0) := (others => '0');5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                          +       v   +    ^	�}     �         2      @    signal rst_count : std_logic(7 downto 0) := (others => '0');5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               $          .       v   .    ^	�     �         2      4    signal rst_count : std_logic := (others => '0');5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                               $          .       v   .    ^	�     �         2      )    signal rst_count : std_logic := '0');5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                               $          .       v   .    ^	�     �         2      (    signal rst_count : std_logic := '0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ^	�   ( �         2                    rst_count <= '1';5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                             ^	�   ) �   #   %   2                     end if;5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^	�   * �   !   #   2      %               --   rst_count <= '0';5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^	�     �   !   #   2      $               -   rst_count <= '0';5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^	�     �   !   #   2      #                  rst_count <= '0';5�_�   �               �   "       ����                                                                                                                                                                                                                                                                                                                                                             ^	��     �   !   #   2      '               iiii   rst_count <= '0';5�_�   [   _   \   `   ^      -    ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	׫     �         .      5                    spi_miso   <= misoSignal(count7);5�_�   ^               _      2    ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	׬    �         .      4                    spi_miso   <= misoSignal(count);5�_�   [   ]       ^   \          ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	��     �         .      K                       internalMmisoSignal <= misoSignal(6 downto 0) & '0';5�_�   \               ]           ����                                                                                                                                                                                                                                                                                                                            (          +          V       ^	��     �         .      J                       internalMisoSignal <= misoSignal(6 downto 0) & '0';5�_�   ,   .       /   -          ����                                                                                                                                                                                                                                                                                                                            +           0                   ^��     �         2      )            else if rising_edge(clk) then5�_�   -               .          ����                                                                                                                                                                                                                                                                                                                            +           0                   ^��     �         1      (            elseif rising_edge(clk) then5��