Vim�UnDo� ���Ac��X�c��.�?�m�ܤ���/�m�   1   end architecture lab1_tb_arq   1         p       p   p   p    ]�=�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                   �               5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                 �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                5�_�      
                      ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                begin5�_�         	       
          ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �               end5�_�   
                    	    ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �               
   end la 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                  end lab1_tb 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �               end lab1_tb 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �   	             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�2     �                  5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�2     �      
            �      
       5�_�                    	        ����                                                                                                                                                                                                                                                                                                                            	           	           V        ]�2-     �             �   	   
       �      	             component 5�_�                    	        ����                                                                                                                                                                                                                                                                                                                            	                     V        ]�2.     �      
   (      entity lab1 is5�_�                            ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2H     �                       begin5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2N     �         &      end entity lab1;5�_�                      .    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2v     �         &      /      led: out std_logic_vector ( 3 downto 0 );5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         �         &    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         signal clk: out5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         signal clk_tb: out5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         signal clk_tb: std_logic_5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         signal clk_tb: std_logic:5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '         signal clk_tb: std_logic:=0;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '          signal clk_tb: std_logic:='0;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         '    �         '    5�_�      !                  
    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         (      !   signal clk_tb: std_logic:='0';5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         )         �         (    5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2�     �         *    �         *    5�_�   "   $           #      
    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�3     �         +      6   signal led_tb: std_logic_vector(3 downto 0):='0000'5�_�   #   %           $           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�3     �                 5�_�   $   &           %   !   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�3B     �       #   *      6         A_tb <= transport vectorA(i) after (tiempo); 5�_�   %   '           &   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�3Y     �   !   #   +    5�_�   &   (           '      4    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�3`     �         ,      6   signal swt_tb: std_logic_vector(3 downto 0):='0000'5�_�   '   )           (   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4_     �       "   ,               swt_tb<='0001'5�_�   (   *           )   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4g     �       "   ,               swt_tb(0)<='0001'5�_�   )   +           *   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4g     �       "   ,               swt_tb(0)<='001'5�_�   *   ,           +   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4h     �       "   ,               swt_tb(0)<='01'5�_�   +   -           ,   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4l     �       "   ,    �   !   "   ,    5�_�   ,   .           -   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4n     �   !   #   -               swt_tb(0)<='1'5�_�   -   /           .   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4o     �   !   #   -               swt_tb(1)<='1'5�_�   .   0           /   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4p     �   !   #   -               swt_tb(1)<=5�_�   /   2           0   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4}     �   !   #   -               swt_tb(1)<=swt_tb(0)l5�_�   0   3   1       2   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �       "   -               swt_tb(0)<='1'5�_�   2   4           3   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �       "   -               swt_tb(0)<='1';5�_�   3   5           4   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   -               swt_tb(1)<=swt_tb(0);5�_�   4   6           5   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   -               swt_tb(3)<=swt_tb(0);5�_�   5   7           6   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   -    �   "   #   -    5�_�   6   8           7   "   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   .    �   "   #   .    5�_�   7   9           8   "   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   /    �   "   #   /    5�_�   8   :           9   "   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   !   #   0    �   "   #   0    5�_�   9   ;           :   #       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   "   $   1               swt_tb(3)<=swt_tb(2);5�_�   :   <           ;   $       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   #   %   1               swt_tb(3)<=swt_tb(2);5�_�   ;   =           <   %       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   $   &   1               swt_tb(3)<=swt_tb(2);5�_�   <   >           =   #       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   "   $   1               swt_tb(2)<=swt_tb(2);5�_�   =   ?           >   $       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   #   %   1               swt_tb(1)<=swt_tb(2);5�_�   >   @           ?   %       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   $   &   1               swt_tb(1)<=swt_tb(2);5�_�   ?   A           @   %       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   $   &   1               swt_tb(1)<=5�_�   @   B           A   &   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �   %   &                   swt_tb(3)<=swt_tb(2);5�_�   A   C           B   !        ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �       !                   swt_tb(3)<='1';5�_�   B   D           C      4    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �         /      6   signal swt_tb: std_logic_vector(3 downto 0):='0001'5�_�   C   E           D      4    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4�     �         /      6   signal swt_tb: std_logic_vector(3 downto 0):='0009'5�_�   D   F           E   %        ����                                                                                                                                                                                                                                                                                                                            %           )   "       V   4    ]�4�     �   $   %           5�_�   E   G           F   $       ����                                                                                                                                                                                                                                                                                                                            %           (   "       V   4    ]�7�     �   $   &   /      	         �   $   &   .    5�_�   F   H           G   &        ����                                                                                                                                                                                                                                                                                                                            &          +          V       ]�7�     �   %   &          >                 A_tb <= transport vectorA(i) after (tiempo);    5         B_tb <= transport vectorB(i) after (tiempo);   1         load_tb <= transport '1' after (tiempo);   "         tiempo := tiempo + 40 ns;   1         load_tb <= transport '0' after (tiempo);   #         tiempo := tiempo + 260 ns;5�_�   G   I           H           ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�    �   (                 end process;�   '   )   )            wait;�   &   (   )            �   %   '   )            end loop;�   $   &   )               wait for 100ns�   #   %   )               swt_tb(1)<='1';�   "   $   )               swt_tb(1)<=swt_tb(0);�   !   #   )               swt_tb(2)<=swt_tb(1);�       "   )               swt_tb(3)<=swt_tb(2);�      !   )            for i in 0 to 6 loop�          )         begin�         )      d      variable vectorB: auxiliar := ("00101", "00001", "00011", "00000", "00100", "01100", "00011");�         )      d      variable vectorA: auxiliar := ("00011", "00010", "01111", "00010", "00000", "01111", "01110");�         )      *      variable tiempo: time      := 15 ns;�         )      
   process�         )         rst_tb <= '0' after 5 ns;�         )      $   clk_tb <= not clk_tb after 25 ns;�         )      6   signal swt_tb: std_logic_vector(3 downto 0):='0000'�         )      6   signal led_tb: std_logic_vector(3 downto 0):='0000'�         )      !   signal rst_tb: std_logic:='0';�         )      !   signal clk_tb: std_logic:='0';�         )         end component lab1;�         )          );�         )      .      led: out std_logic_vector ( 3 downto 0 )�         )      /      swt: in  std_logic_vector ( 3 downto 0 );�         )      	   port (�         )         );�   
      )         N:=1�   	      )         generic (�      
   )         component lab1 is�                %      variable tiempo: time := 15 ns;�                d      variable vectorB: auxiliar := ("00101", "00001", "00011", "00000", "00100", "01100", "00011");�                d      variable vectorA: auxiliar := ("00011", "00010", "01111", "00010", "00000", "01111", "01110");5�_�   H   K           I   '        ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   &   (   )            5�_�   I   L   J       K   '        ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   &   '           5�_�   K   M           L   '       ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   &   (   (            wait;5�_�   L   N           M   (       ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   (            �   (            5�_�   M   O           N   )        ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   (               5�_�   N   Q           O   )       ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�    �   (              end entity lab1_tb_arq5�_�   O   R   P       Q           ����                                                                                                                                                                                                                                                                                                                                                  V        ]�<     �                *      variable tiempo: time      := 15 ns;   d      variable vectorA: auxiliar := ("00011", "00010", "01111", "00010", "00000", "01111", "01110");   d      variable vectorB: auxiliar := ("00101", "00001", "00011", "00000", "00100", "01100", "00011");5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                                                             ]�<r     �         &    �         &    5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                                                             ]�<v     �                library ieee;5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                                                             ]�<w     �                use ieee.std_logic_1164.all;5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                             ]�<y    �         '      use IEEE.std_logic_1164.all.5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                             ]�<�     �         '         end component lab1;5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                             ]�<�     �         '         end component ;5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                                                             ]�<�     �         '         N:=15�_�   X   Z           Y   &       ����                                                                                                                                                                                                                                                                                                                                                             ]�<�     �   %   )   '         end process;5�_�   Y   [           Z   (       ����                                                                                                                                                                                                                                                                                                                                                             ]�=     �   '   )   )         aaa:lab1_tb5�_�   Z   \           [   (       ����                                                                                                                                                                                                                                                                                                                                                             ]�=     �   '   *   )         aaa:lab15�_�   [   ]           \   )       ����                                                                                                                                                                                                                                                                                                                                                             ]�=     �   (   *   *         map5�_�   \   ^           ]   )   	    ����                                                                                                                                                                                                                                                                                                                                                             ]�=     �   (   *   *         generica map5�_�   ]   _           ^   )   	    ����                                                                                                                                                                                                                                                                                                                                                             ]�=      �   (   *   *         generia map5�_�   ^   `           _   )       ����                                                                                                                                                                                                                                                                                                                                                             ]�=$     �   (   ,   *         generic map5�_�   _   a           `   *       ����                                                                                                                                                                                                                                                                                                                                                             ]�=3     �   )   +   ,            N => 4;5�_�   `   b           a   +        ����                                                                                                                                                                                                                                                                                                                                                             ]�=4     �   *   ,          );5�_�   a   c           b   +       ����                                                                                                                                                                                                                                                                                                                                                             ]�=9     �   +   .   -         �   +   -   ,    5�_�   b   d           c   -        ����                                                                                                                                                                                                                                                                                                                                                V       ]�=I     �   ,   /   .    �   -   .   .    5�_�   c   e           d   -   	    ����                                                                                                                                                                                                                                                                                                                            -   	       .   	          	    ]�=M     �   -   /   0      .      led: out std_logic_vector ( 3 downto 0 )�   ,   .   0      /      swt: in  std_logic_vector ( 3 downto 0 );5�_�   d   f           e   -   	    ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=V     �   ,   .   0      /      swt: in  std_logic_vector ( 3 downto 0 );�   ,   /   0      1      swt<=: in  std_logic_vector ( 3 downto 0 );   0      led<=: out std_logic_vector ( 3 downto 0 )5�_�   e   g           f   -       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=]     �   ,   .   0      1      swt=>: in  std_logic_vector ( 3 downto 0 );5�_�   f   h           g   -       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=c     �   ,   .   0      7      swt=>swt_tb: in  std_logic_vector ( 3 downto 0 );5�_�   g   i           h   .       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=e     �   -   /   0      0      led=>: out std_logic_vector ( 3 downto 0 )5�_�   h   j           i   .       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=j     �   -   /   0      6      led=>led_tb: out std_logic_vector ( 3 downto 0 )5�_�   i   k           j   -       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=o     �   ,   .   0      7      swt=>swt_tb; in  std_logic_vector ( 3 downto 0 );5�_�   j   l           k   .       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=p     �   -   /   0      6      led=>led_tb; out std_logic_vector ( 3 downto 0 )5�_�   k   m           l   -       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=q     �   ,   .   0      7      swt=>swt_tb, in  std_logic_vector ( 3 downto 0 );5�_�   l   n           m   .       ����                                                                                                                                                                                                                                                                                                                            -   	       .   
          
    ]�=r     �   .   0   1            �   .   0   0    5�_�   m   o           n   *        ����                                                                                                                                                                                                                                                                                                                            )          /          V       ]�=�     �   .   0             )r�   -   /                led=>led_tb�   ,   .                swt=>swt_tb,�   *   ,             );�   )   +                N => 45�_�   n   p           o   /       ����                                                                                                                                                                                                                                                                                                                            )          /          V       ]�=�     �   .   0   1                  )r5�_�   o               p   1       ����                                                                                                                                                                                                                                                                                                                            )          /          V       ]�=�    �   0              end architecture lab1_tb_arq5�_�   O           Q   P      
    ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �         )         process myProcces5�_�   I           K   J   (        ����                                                                                                                                                                                                                                                                                                                                                V       ]�7�     �   '   )        5�_�   0           2   1   !       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�4~     �       "   -               swt_tb(0)<='1;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�2o     �         &            5�_�              
   	          ����                                                                                                                                                                                                                                                                                                                                                             ]�1�     �                  end 5��