Vim�UnDo� �
Lm�T�su��A�a�նӒ�C�~����   =   )           n_axis_tready : in  STD_LOGIC;            �       �   �   �    ^�    _�                            ����                                                                                                                                                                                                                                                                                                                                                             ^˶     �         @      entity stretcher is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^˾     �         @      end stretcher;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ^��    �         @      'architecture Behavioral of stretcher is5�_�                    -        ����                                                                                                                                                                                                                                                                                                                            -          :          V       ^��     �   ,   ;   @    �   -   .   @    5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            ;          H          V       ^��     �   ,   .   N      $               when waitingMready =>5�_�                    /       ����                                                                                                                                                                                                                                                                                                                            /          /   !       v   !    ^Ӥ     �   .   0   N      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   /   0   N    5�_�                    *   &    ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^Ӿ     �   )   +   N      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�      	              1       ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^��     �   0   1          t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�      
           	   1   %    ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^��     �   0   2   M      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�   	              
   1   /    ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^�      �   0   2   M      b                        m_axis_tdata(bitCounter0) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�   
                 1   A    ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^�     �   0   2   M      a                        m_axis_tdata(bitCounter) <= s_axis_tdata(bitCounter);    --pongo el dato 5�_�                    1   A    ����                                                                                                                                                                                                                                                                                                                            )          )   !       v   !    ^�     �   0   2   M      X                        m_axis_tdata(bitCounter) <= s_axis_tdata(1);    --pongo el dato 5�_�                   1        ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�     �   J   L   M         end process shift_reg;�   I   K   M            end if;�   H   J   M               end if;�   G   I   M                  end case;�   F   H   M                        end if;�   E   G   M      �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   D   F   M                        else�   C   E   M                           end if;�   B   D   M      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar�   A   C   M      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   @   B   M                           else�   ?   A   M      T                        bitCounter      := bitCounter+1;                --incremento�   >   @   M      X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato �   =   ?   M      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   <   >   M      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   ;   =   M      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   :   <   M      }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   9   ;   M      $               when waitingMready =>�   8   :   M                        end if;�   7   9   M      �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)�   6   8   M                        else�   5   7   M                           end if;�   4   6   M      r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar�   3   5   M      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   2   4   M                           else�   1   3   M      ]                        bitCounter               := bitCounter+1;                --incremento�   0   2   M      S                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);--pongo el dato�   /   1   M      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   .   0   M      q                  if s_axis_tvalid = '1' then                           --lo puedo empezar a mandar al otro lado?�   -   /   M      }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora�   ,   .   M      "               when readingData =>�   +   -   M                        end if;�   *   ,   M      (                     bitCounter    := 0;�   )   +   M      �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato�   (   *   M      i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo�   '   )   M      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   M      $               when waitingSvalid =>�   %   '   M                  case state is�   $   &   M               else�   #   %   M      -            m_axis_tdata  <= (others => '0');�   "   $   M      !            m_axis_tvalid <= '0';�   !   #   M      !            s_axis_tready <= '0';�       "   M      +            state         <= waitingSvalid;�      !   M               if rst = '0' then�          M            if rising_edge(clk) then�         M         begin�         M      0      variable bitCounter :integer range 0 to 8;�         M         shift_reg:process (clk) is�         M      ,   signal state:shiftState := waitingSvalid;�         M      5   type shiftState is (waitingSvalid, waitingMready);�         M      *           rst           : in  STD_LOGIC);�         M      )           clk           : in  STD_LOGIC;�         M      )           s_axis_tready : out STD_LOGIC;�         M      )           s_axis_tlast  : in  STD_LOGIC;�         M      )           s_axis_tvalid : in  STD_LOGIC;�         M      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         M      )           m_axis_tready : in  STD_LOGIC;�   
      M      )           m_axis_tlast  : out STD_LOGIC;�   	      M      )           m_axis_tvalid : out STD_LOGIC;�      
   M      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   M          Port(  �   0   2          X                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);    --pongo el dato �   1   3          T                        bitCounter      := bitCounter+1;                --incremento5�_�                    1   D    ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�      �   0   2   M      S                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);--pongo el dato5�_�                    2   G    ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�#     �   1   3   M      ]                        bitCounter               := bitCounter+1;                --incremento5�_�                   2   G    ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�'     �   1   3   M      S                        bitCounter               := bitCounter+1;      --incremento5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�4     �   -   .          }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�                    6        ����                                                                                                                                                                                                                                                                                                                            6          7          V       ^�O     �   5   6                            else   �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)5�_�                    3   0    ����                                                                                                                                                                                                                                                                                                                            6          6          V       ^�b     �   2   4   J      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�                    3   1    ����                                                                                                                                                                                                                                                                                                                            6          6          V       ^�e     �   2   4   J      m                        state         <= waitingMvalid;                 --termine de mandar, vuelvo a esperar5�_�                    3   6    ����                                                                                                                                                                                                                                                                                                                            6          6          V       ^�f     �   2   4   J      r                        state         <= waitingMreadyvalid;                 --termine de mandar, vuelvo a esperar5�_�                    4        ����                                                                                                                                                                                                                                                                                                                            4          4          V       ^�p     �   3   5   I    �   4   5   I    �   3   4          r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            4           4   h       V       ^�q     �   3   5   J      i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�                    4   *    ����                                                                                                                                                                                                                                                                                                                            4           4   h       V       ^ض     �   3   5   J      l                        s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�                    4   *    ����                                                                                                                                                                                                                                                                                                                            4           4   h       V       ^��     �   3   5   J    �   4   5   J    5�_�                    5       ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   4   6   K      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�                    5       ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   4   6   K      l                        m_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�                     5        ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   4   6   K      l                        m_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�      !               5   *    ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   4   6   K      l                        m_axis_tvalid <= '0';                              --entonces yo tambien estoy listo5�_�       "           !   5   -    ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   4   6   K      l                        m_axis_tvalid <= '1';                              --entonces yo tambien estoy listo5�_�   !   #           "   4   -    ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   3   5   K      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�   "   $           #   3   7    ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   2   4   K      m                        state         <= waitingMready;                 --termine de mandar, vuelvo a esperar5�_�   #   %           $   9       ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   8   9          }                     s_axis_tready <= '0';                              --el dato esta en la mesa, ya no quiero mas por ahora5�_�   $   &           %   :       ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   9   ;   J    �   :   ;   J    5�_�   %   '           &   :   *    ����                                                                                                                                                                                                                                                                                                                            5           5   h       V       ^��     �   9   ;   K      -                        m_axis_tvalid <= '1';5�_�   &   (           '   ;        ����                                                                                                                                                                                                                                                                                                                            ;          ?          V       ^��     �   :   ;          f                     if bitCounter < 8 then                             --perfecto, porque bit voy?      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato   X                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato    T                        bitCounter      := bitCounter+1;                --incremento                        else5�_�   '   )           (   <       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^��     �   ;   <          r                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar5�_�   (   *           )   <       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^�      �   ;   <                               end if;5�_�   )   ,           *   <        ����                                                                                                                                                                                                                                                                                                                            <          =          V       ^�    �   ;   <                            else   �                     m_axis_tvalid <= '0';                              --si en la mitad de la transmision el receptor no puede recibir, lo espero (pero me ofendo y yo tampoco transmito)5�_�   *   -   +       ,      &    ����                                                                                                                                                                                                                                                                                                                            <          <          V       ^�     �         B      5   type shiftState is (waitingSvalid, waitingMready);�         B    5�_�   ,   /           -      1    ����                                                                                                                                                                                                                                                                                                                            <          <          V       ^��    �         B      @   type shiftState is (waitingSvalid, readingDatawaitingMready);5�_�   -   0   .       /          ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �         B      I--tomo 1 byte y mando 8 bytes en donde en cada uno de salida vale el bit05�_�   /   1           0      W    ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �         B      �--junto 8 bytes en uno, tomando solo el bit 0 de cada byte y lo mando por el axi mastertomo 1 byte y mando 8 bytes en donde en cada uno de salida vale el bit05�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �                ?-- lo hago para entrar al convolucionador que recibe de a 1 but5�_�   1   3           2   -   J    ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �   ,   .   A      q                  if s_axis_tvalid = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�   2   4           3   -   J    ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �   ,   .   A      J                  if s_axis_tvalid = '1' then                           --5�_�   3   5           4   .   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�     �   -   /   A      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�   4   6           5   /   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�     �   .   0   A      W                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);    --pongo el dato5�_�   5   7           6   /   g    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�     �   .   0   A      t                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);    --voy armando el dato but a butpongo el dato5�_�   6   8           7   2   7    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�"     �   1   3   A      7                        state         <= waitingMready;5�_�   7   9           8   3   -    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�,     �   2   4   A      -                        s_axis_tready <= '0';5�_�   8   :           9   4   -    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�:     �   3   5   A      -                        m_axis_tvalid <= '1';5�_�   9   ;           :   8   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�G     �   7   9   A      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�   :   <           ;   8   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�G     �   7   9   A      J                  if m_axis_tready = '1' then                           --5�_�   ;   =           <   9   -    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�R     �   8   :   A      -                        m_axis_tvalid <= '0';5�_�   <   >           =   8   f    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�X     �   7   9   A      h                  if m_axis_tready = '1' then                           --si el receptor puede recibir..5�_�   =   ?           >   9   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�c     �   8   :   A      J                        m_axis_tvalid <= '0';                           --5�_�   >   @           ?   :   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�j     �   9   ;   A      m                        state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�   ?   A           @   :   J    ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^�k    �   9   ;   A      J                        state         <= waitingSvalid;                 --5�_�   @   B           A   !       ����                                                                                                                                                                                                                                                                                                                            .   J       .   S       v   S    ^��     �       "   A      !            s_axis_tready <= '0';5�_�   A   C           B   (        ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   '   (          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   B   D           C   9       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   8   :   @    �   9   :   @    5�_�   C   E           D   9       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   8   :          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   D   F           E   9   G    ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   8   :   A      l                        s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   E   G           F   9   I    ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   8   :   A      h                        s_axis_tready <= '1';                          --entonces yo tambien estoy listo5�_�   F   H           G   9   G    ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��    �   8   :   A      i                        s_axis_tready <= '1';                          -- entonces yo tambien estoy listo5�_�   G   I           H   .   %    ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^�    �   -   /   A      g                        m_axis_tdata(bitCounter) <= s_axis_tdata(0);    --voy armando el dato but a but5�_�   H   J           I   $        ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^�{     �   #   %   A    �   $   %   A    5�_�   I   K           J   $       ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�|     �   #   %          (                     bitCounter    := 0;5�_�   J   L           K   ;   (    ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�     �   :   <   B      Z                        state         <= waitingSvalid;                 --cambio de estado5�_�   K   M           L   ;   5    ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�     �   :   <   B      W                        state         <=readingData;                 --cambio de estado5�_�   L   N           M   ;   8    ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�     �   :   <   B      [                        state         <=readingData;                     --cambio de estado5�_�   M   O           N   &        ����                                                                                                                                                                                                                                                                                                                            &          +          V   )    ^�     �   %   &                      case state is   $               when waitingSvalid =>   r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato   (                     bitCounter    := 0;                     end if;5�_�   N   P           O           ����                                                                                                                                                                                                                                                                                                                            &          &          V   )    ^�     �      !   <      +            state         <= waitingSvalid;5�_�   O   Q           P   )        ����                                                                                                                                                                                                                                                                                                                            )   '       *   '       V   '    ^�     �   9   ;   <         end process shift_reg;�   8   :   <            end if;�   7   9   <               end if;�   6   8   <                  end case;�   5   7   <                        end if;�   4   6   <      Z                        state         <=readingData;                    --cambio de estado�   3   5   <      j                        s_axis_tready <= '1';                           -- entonces yo tambien estoy listo�   2   4   <      `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   1   3   <      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   0   2   <      $               when waitingMready =>�   /   1   <                        end if;�   .   0   <                           end if;�   -   /   <      b                        m_axis_tvalid <= '1';                           -- pero si para transmitir�   ,   .   <      o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos�   +   -   <      d                        state         <= waitingMready;                 -- termine, cambio de estado�   *   ,   <                           else�   )   +   <      V                        bitCounter                 := bitCounter+1;       --incremento�   (   *   <      e                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);--voy armando el dato but a but�   '   )   <      \                     if bitCounter < 8 then                             --porque bit voy?   �   &   (   <      u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte�   %   '   <      "               when readingData =>�   $   &   <               else�   #   %   <                  bitCounter    := 0;�   "   $   <      -            m_axis_tdata  <= (others => '0');�   !   #   <      !            m_axis_tvalid <= '0';�       "   <      !            s_axis_tready <= '1';�      !   <      )            state         <= readingData;�          <               if rst = '0' then�         <            if rising_edge(clk) then�         <         begin�         <      0      variable bitCounter :integer range 0 to 8;�         <         shift_reg:process (clk) is�         <      ,   signal state:shiftState := waitingSvalid;�         <      B   type shiftState is (waitingSvalid, readingData, waitingMready);�         <      *           rst           : in  STD_LOGIC);�         <      )           clk           : in  STD_LOGIC;�         <      )           s_axis_tready : out STD_LOGIC;�         <      )           s_axis_tlast  : in  STD_LOGIC;�         <      )           s_axis_tvalid : in  STD_LOGIC;�         <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      <      )           m_axis_tready : in  STD_LOGIC;�   	      <      )           m_axis_tlast  : out STD_LOGIC;�      
   <      )           m_axis_tvalid : out STD_LOGIC;�      	   <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         <          Port(  �   (   *          i                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);    --voy armando el dato but a but�   )   +          T                        bitCounter               := bitCounter+1;       --incremento5�_�   P   R           Q   )   F    ����                                                                                                                                                                                                                                                                                                                            )   '       *   '       V   '    ^�     �   (   *   <      e                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);--voy armando el dato but a but5�_�   Q   S           R   *   G    ����                                                                                                                                                                                                                                                                                                                            )   '       *   '       V   '    ^�     �   )   +   <      V                        bitCounter                 := bitCounter+1;       --incremento5�_�   R   T           S   *   G    ����                                                                                                                                                                                                                                                                                                                            )   '       *   '       V   '    ^�    �   )   +   <      U                        bitCounter                 := bitCounter+1;      --incremento5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ^��     �         <      B   type shiftState is (waitingSvalid, readingData, waitingMready);5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ^��   	 �         <      ,   signal state:shiftState := waitingSvalid;5�_�   U   W           V   5       ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ^��     �   4   6   <    �   5   6   <    5�_�   V   X           W   5       ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ^��     �   4   6                      bitCounter    := 0;5�_�   W   Y           X   3        ����                                                                                                                                                                                                                                                                                                                            3          6          V       ^��     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      [                        state         <= readingData;                    --cambio de estado�   4   6   =      +                        bitCounter    := 0;�   3   5   =      j                        s_axis_tready <= '1';                           -- entonces yo tambien estoy listo�   2   4   =      E                        m_axis_tvalid <= '0';--y ya no tengo mas nada�   1   3   =      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   0   2   =      $               when waitingMready =>�   /   1   =                        end if;�   .   0   =                           end if;�   -   /   =      b                        m_axis_tvalid <= '1';                           -- pero si para transmitir�   ,   .   =      o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos�   +   -   =      d                        state         <= waitingMready;                 -- termine, cambio de estado�   *   ,   =                           else�   )   +   =      T                        bitCounter                 := bitCounter+1;     --incremento�   (   *   =      g                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);  --voy armando el dato but a but�   '   )   =      \                     if bitCounter < 8 then                             --porque bit voy?   �   &   (   =      u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte�   %   '   =      "               when readingData =>�   $   &   =               else�   #   %   =                  bitCounter    := 0;�   "   $   =      -            m_axis_tdata  <= (others => '0');�   !   #   =      !            m_axis_tvalid <= '0';�       "   =      !            s_axis_tready <= '1';�      !   =      )            state         <= readingData;�          =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      *   signal state:shiftState := readingData;�         =      3   type shiftState is (readingData, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      =      )           m_axis_tready : in  STD_LOGIC;�   	      =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   2   4          `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   5   7          Z                        state         <=readingData;                    --cambio de estado�   4   6          +                        bitCounter    := 0;�   3   5          j                        s_axis_tready <= '1';                           -- entonces yo tambien estoy listo5�_�   X   Z           Y   3   -    ����                                                                                                                                                                                                                                                                                                                            3          6          V       ^��   
 �   2   4   =      E                        m_axis_tvalid <= '0';--y ya no tengo mas nada5�_�   Y   [           Z   &        ����                                                                                                                                                                                                                                                                                                                            3          6          V       ^�,    �   %   '   =    �   &   '   =    5�_�   Z   \           [   )   %    ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�5     �   (   *   >      \                     if bitCounter < 8 then                             --porque bit voy?   5�_�   [   ]           \   )   %    ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�A     �   (   *   >      \                     if bitCounter < 7 then                             --porque bit voy?   5�_�   \   ^           ]   +   %    ����                                                                                                                                                                                                                                                                                                                            4          7          V       ^�C     �   +   .   ?                              �   +   -   >    5�_�   ]   _           ^   ,   (    ����                                                                                                                                                                                                                                                                                                                            6          9          V       ^�l     �   +   -   @      .                        if bitCounter = 8 then5�_�   ^   `           _   ,   (    ����                                                                                                                                                                                                                                                                                                                            6          9          V       ^�p     �   +   -   @      .                        if bitCounter = 8 then5�_�   _   a           `   ,   (    ����                                                                                                                                                                                                                                                                                                                            6          9          V       ^�s     �   ,   .   @    5�_�   `   b           a   -        ����                                                                                                                                                                                                                                                                                                                            7          :          V       ^�y     �   -   /   A    �   -   .   A    5�_�   a   c           b   -        ����                                                                                                                                                                                                                                                                                                                            8          ;          V       ^�z     �   ,   -           5�_�   b   d           c   -       ����                                                                                                                                                                                                                                                                                                                            7          :          V       ^�{     �   ,   .          o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos5�_�   c   e           d   .        ����                                                                                                                                                                                                                                                                                                                            7          :          V       ^�|     �   -   .           5�_�   d   f           e   !       ����                                                                                                                                                                                                                                                                                                                            6          9          V       ^�     �       "   @      !            s_axis_tready <= '1';5�_�   e   g           f   '        ����                                                                                                                                                                                                                                                                                                                            '          3          V       ^�5     �   &   4   @    �   '   (   @    5�_�   f   h           g   '        ����                                                                                                                                                                                                                                                                                                                            '           3           V        ^�?     �   &   -   @    �   '   (   @    �   &   '          "               when readingData =>   u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte   \                     if bitCounter < 8 then                             --porque bit voy?      g                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);  --voy armando el dato but a but   T                        bitCounter                 := bitCounter+1;     --incremento   .                        if bitCounter = 7 then   r                           s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos                        else   d                        state         <= waitingMready;                 -- termine, cambio de estado   o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos   b                        m_axis_tvalid <= '1';                           -- pero si para transmitir                        end if;                     end if;5�_�   g   i           h   *   &    ����                                                                                                                                                                                                                                                                                                                            '           ,          V        ^��     �   )   +   F      �                     state         <= waitingMready;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   h   j           i   $       ����                                                                                                                                                                                                                                                                                                                            '           ,          V        ^��     �   #   $                      bitCounter    := 0;5�_�   i   k           j           ����                                                                                                                                                                                                                                                                                                                            &           +          V        ^��     �      !   E      )            state         <= readingData;5�_�   j   l           k   1        ����                                                                                                                                                                                                                                                                                                                            1   %       2   %       V   %    ^��     �   0   1          .                        if bitCounter = 7 then   r                           s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos5�_�   k   m           l   :       ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �   9   :          j                        s_axis_tready <= '1';                           -- entonces yo tambien estoy listo5�_�   l   n           m   :       ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �   9   :          +                        bitCounter    := 0;5�_�   m   o           n   :   )    ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �   9   ;   A      [                        state         <= readingData;                    --cambio de estado5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��     �         A      3   type shiftState is (readingData, waitingMready);5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                            1   %       1   %       V   %    ^��    �         A      *   signal state:shiftState := readingData;5�_�   p   s           q   /        ����                                                                                                                                                                                                                                                                                                                            /           0           V        ^ �     �   .   1   A      g                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);  --voy armando el dato but a but   T                        bitCounter                 := bitCounter+1;     --incremento5�_�   q   t   r       s   (        ����                                                                                                                                                                                                                                                                                                                            /           0           V        ^ �     �   '   *   A    �   (   )   A    5�_�   s   u           t   (        ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^ �     �   (   *          T                        bitcounter                 := bitcounter+1;     --incremento�   '   )          g                        m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);  --voy armando el dato but a but5�_�   t   v           u   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^ �     �   +   ,          (                     bitCounter    := 0;5�_�   u   w           v   (       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^ �     �   '   )   B    �   (   )   B    5�_�   v   x           w   *   "    ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^;     �   )   +   C    �   *   +   C    5�_�   w   y           x   )        ����                                                                                                                                                                                                                                                                                                                            *          )          V       ^>     �   A   C   D         end process shift_reg;�   @   B   D            end if;�   ?   A   D               end if;�   >   @   D                  end case;�   =   ?   D                        end if;�   <   >   D      ]                        state         <= waitingSvalid;                    --cambio de estado�   ;   =   D      `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   :   <   D      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   9   ;   D      $               when waitingMready =>�   8   :   D                        end if;�   7   9   D                           end if;�   6   8   D      b                        m_axis_tvalid <= '1';                           -- pero si para transmitir�   5   7   D      o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos�   4   6   D      d                        state         <= waitingMready;                 -- termine, cambio de estado�   3   5   D                           else�   2   4   D      T                        bitcounter                 := bitcounter+1;     --incremento�   1   3   D      g                        m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);  --voy armando el dato but a but�   0   2   D      \                     if bitCounter < 8 then                             --porque bit voy?   �   /   1   D      u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte�   .   0   D      "               when readingData =>�   -   /   D                        end if;�   ,   .   D      �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato�   +   -   D      i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo�   *   ,   D      Q                     bitcounter                 := bitcounter+1;     --incremento�   )   +   D      i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo�   (   *   D      b                     m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);--voy armando el dato but a but�   '   )   D      (                     bitCounter    := 0;�   &   (   D      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   %   '   D      $               when waitingSvalid =>�   $   &   D                  case state is�   #   %   D               else�   "   $   D      -            m_axis_tdata  <= (others => '0');�   !   #   D      !            m_axis_tvalid <= '0';�       "   D      !            s_axis_tready <= '0';�      !   D      +            state         <= waitingSvalid;�          D               if rst = '0' then�         D            if rising_edge(clk) then�         D         begin�         D      0      variable bitCounter :integer range 0 to 8;�         D         shift_reg:process (clk) is�         D      ,   signal state:shiftState := waitingSvalid;�         D      B   type shiftState is (waitingSvalid, readingData, waitingMready);�         D      *           rst           : in  STD_LOGIC);�         D      )           clk           : in  STD_LOGIC;�         D      )           s_axis_tready : out STD_LOGIC;�         D      )           s_axis_tlast  : in  STD_LOGIC;�         D      )           s_axis_tvalid : in  STD_LOGIC;�         D      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      D      )           m_axis_tready : in  STD_LOGIC;�   	      D      )           m_axis_tlast  : out STD_LOGIC;�      
   D      )           m_axis_tvalid : out STD_LOGIC;�      	   D      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         D          Port(  �   (   *          d                     m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);  --voy armando el dato but a but5�_�   x   z           y   )   C    ����                                                                                                                                                                                                                                                                                                                            *          )          V       ^A     �   (   *   D      b                     m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);--voy armando el dato but a but5�_�   y   {           z   +       ����                                                                                                                                                                                                                                                                                                                            *          )          V       ^F     �   *   +          Q                     bitcounter                 := bitcounter+1;     --incremento5�_�   z   |           {   +       ����                                                                                                                                                                                                                                                                                                                            *          )          V       ^I     �   *   +          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   {   }           |   (       ����                                                                                                                                                                                                                                                                                                                            *          )          V       ^d     �   '   (          (                     bitCounter    := 0;5�_�   |   ~           }   )       ����                                                                                                                                                                                                                                                                                                                            )          (          V       ^r     �   (   *   A    �   )   *   A    5�_�   }              ~   (       ����                                                                                                                                                                                                                                                                                                                            *          (          V       ^�     �   (   *   B    �   (   )   B    5�_�   ~   �              )       ����                                                                                                                                                                                                                                                                                                                            +          (          V       ^�     �   (   *   C      \                     if bitCounter < 8 then                             --porque bit voy?   5�_�      �           �   )       ����                                                                                                                                                                                                                                                                                                                            +          (          V       ^�     �   (   *   C                           5�_�   �   �           �   (   '    ����                                                                                                                                                                                                                                                                                                                            +          (          V       ^�     �   '   )   C      C                     m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            +          (          V       ^�     �   (   *   C                           bitCounter5�_�   �   �           �   )   1    ����                                                                                                                                                                                                                                                                                                                            +          (          V       ^�     �   (   *   C      2                     bitCounter := bitCounter + 1:5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�     �   *   +          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�     �   (   *   B    �   )   *   B    5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�     �   '   )   C    �   (   )   C    5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^�     �   )   +          i                     s_axis_tready <= '1';                              --entonces yo tambien estoy listo�   (   *          C                     m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   *   '    ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^     �   *   ,   E                              �   *   ,   D    5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^/     �   +   -   E    �   ,   -   E    5�_�   �   �           �   ,   *    ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^1     �   +   -   F      l                        s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /   *       /   *       V   *    ^?     �   .   /          �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            /   *       /   *       V   *    ^?     �   ,   .   E    �   -   .   E    5�_�   �   �   �       �   +       ����                                                                                                                                                                                                                                                                                                                            0   *       0   *       V   *    ^T     �   *   ,   F    �   +   ,   F    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            1   *       1   *       V   *    ^U     �   *   ,          2                     bitCounter := bitCounter + 1;5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^X     �   D   F   G         end process shift_reg;�   C   E   G            end if;�   B   D   G               end if;�   A   C   G                  end case;�   @   B   G                        end if;�   ?   A   G      ]                        state         <= waitingSvalid;                    --cambio de estado�   >   @   G      `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   =   ?   G      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   <   >   G      $               when waitingMready =>�   ;   =   G                        end if;�   :   <   G                           end if;�   9   ;   G      b                        m_axis_tvalid <= '1';                           -- pero si para transmitir�   8   :   G      o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos�   7   9   G      d                        state         <= waitingMready;                 -- termine, cambio de estado�   6   8   G                           else�   5   7   G      T                        bitcounter                 := bitcounter+1;     --incremento�   4   6   G      g                        m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);  --voy armando el dato but a but�   3   5   G      \                     if bitCounter < 8 then                             --porque bit voy?   �   2   4   G      u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte�   1   3   G      "               when readingData =>�   0   2   G                        end if;�   /   1   G      \                     if bitCounter < 8 then                             --porque bit voy?   �   .   0   G      2                     bitCounter := bitCounter + 1;�   -   /   G      �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato�   ,   .   G      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   +   -   G                           else �   *   ,   G      E                        bitCounter                 := bitCounter + 1;�   )   +   G      y                        s_axis_tready              <= '1';                              --entonces yo tambien estoy listo�   (   *   G      F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);�   '   )   G      \                     if bitCounter < 8 then                             --porque bit voy?   �   &   (   G      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   %   '   G      $               when waitingSvalid =>�   $   &   G                  case state is�   #   %   G               else�   "   $   G      -            m_axis_tdata  <= (others => '0');�   !   #   G      !            m_axis_tvalid <= '0';�       "   G      !            s_axis_tready <= '0';�      !   G      +            state         <= waitingSvalid;�          G               if rst = '0' then�         G            if rising_edge(clk) then�         G         begin�         G      0      variable bitCounter :integer range 0 to 8;�         G         shift_reg:process (clk) is�         G      ,   signal state:shiftState := waitingSvalid;�         G      B   type shiftState is (waitingSvalid, readingData, waitingMready);�         G      *           rst           : in  STD_LOGIC);�         G      )           clk           : in  STD_LOGIC;�         G      )           s_axis_tready : out STD_LOGIC;�         G      )           s_axis_tlast  : in  STD_LOGIC;�         G      )           s_axis_tvalid : in  STD_LOGIC;�         G      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      G      )           m_axis_tready : in  STD_LOGIC;�   	      G      )           m_axis_tlast  : out STD_LOGIC;�      
   G      )           m_axis_tvalid : out STD_LOGIC;�      	   G      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         G          Port(  �   (   *          F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);�   *   ,          5                        bitCounter := bitCounter + 1;�   )   +          l                        s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^a     �   .   /          2                     bitCounter := bitCounter + 1;5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   -   /          �                     state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   .   /          \                     if bitCounter < 8 then                             --porque bit voy?   5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   .   0   E    �   /   0   E    5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   .   0                            end if;5�_�   �   �           �   .   )    ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   -   /   F      �                        state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �   .   )    ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   -   /   F      y                        state         <= D;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �   .   )    ����                                                                                                                                                                                                                                                                                                                            +          )          V       ^�     �   -   /   F      )                        state         <= 5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            1          ;          V       ^�     �   0   1          "               when readingData =>   u                  if s_axis_tvalid = '1' then                           --si sigue listo, entonces puedo leer un byte   \                     if bitCounter < 8 then                             --porque bit voy?      g                        m_axis_tdata(7-bitcounter) <= s_axis_tdata(0);  --voy armando el dato but a but   T                        bitcounter                 := bitcounter+1;     --incremento                        else   d                        state         <= waitingMready;                 -- termine, cambio de estado   o                        s_axis_tready <= '0';                           -- ya no estoy listo para recibir datos   b                        m_axis_tvalid <= '1';                           -- pero si para transmitir                        end if;                     end if;5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ^�     �   -   /   ;    �   .   /   ;    5�_�   �   �           �   .   *    ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^�     �   -   /   <      `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada5�_�   �   �           �   5   &    ����                                                                                                                                                                                                                                                                                                                            2          2          V       ^�     �   5   7   =                              �   5   7   <    5�_�   �   �           �   5        ����                                                                                                                                                                                                                                                                                                                            6   '       5   '       V   '    ^�     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      (                        bitCounter := 0;�   4   6   =      F                        state      <= waitingSvalid;--cambio de estado�   3   5   =      `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   2   4   =      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   1   3   =      $               when waitingMready =>�   0   2   =                        end if;�   /   1   =                           end if;�   .   0   =      7                        state         <= waitingMready;�   -   /   =      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   ,   .   =      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   +   -   =                           else �   *   ,   =      E                        bitCounter                 := bitCounter + 1;�   )   +   =      y                        s_axis_tready              <= '1';                              --entonces yo tambien estoy listo�   (   *   =      F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);�   '   )   =      \                     if bitCounter < 8 then                             --porque bit voy?   �   &   (   =      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   %   '   =      $               when waitingSvalid =>�   $   &   =                  case state is�   #   %   =               else�   "   $   =      -            m_axis_tdata  <= (others => '0');�   !   #   =      !            m_axis_tvalid <= '0';�       "   =      !            s_axis_tready <= '0';�      !   =      +            state         <= waitingSvalid;�          =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      B   type shiftState is (waitingSvalid, readingData, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      =      )           m_axis_tready : in  STD_LOGIC;�   	      =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   4   6          ]                        state         <= waitingSvalid;                    --cambio de estado�   5   7          (                        bitCounter := 0;5�_�   �   �           �   5   4    ����                                                                                                                                                                                                                                                                                                                            6   '       5   '       V   '    ^�     �   4   6   =      F                        state      <= waitingSvalid;--cambio de estado5�_�   �   �           �   4        ����                                                                                                                                                                                                                                                                                                                            4   3       6   (       V   3    ^�     �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      +                        bitCounter    := 0;�   4   6   =      7                        state         <= waitingSvalid;�   3   5   =      E                        m_axis_tvalid <= '0';--y ya no tengo mas nada�   2   4   =      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   1   3   =      $               when waitingMready =>�   0   2   =                        end if;�   /   1   =                           end if;�   .   0   =      7                        state         <= waitingMready;�   -   /   =      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   ,   .   =      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   +   -   =                           else �   *   ,   =      E                        bitCounter                 := bitCounter + 1;�   )   +   =      y                        s_axis_tready              <= '1';                              --entonces yo tambien estoy listo�   (   *   =      F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);�   '   )   =      \                     if bitCounter < 8 then                             --porque bit voy?   �   &   (   =      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   %   '   =      $               when waitingSvalid =>�   $   &   =                  case state is�   #   %   =               else�   "   $   =      -            m_axis_tdata  <= (others => '0');�   !   #   =      !            m_axis_tvalid <= '0';�       "   =      !            s_axis_tready <= '0';�      !   =      +            state         <= waitingSvalid;�          =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      B   type shiftState is (waitingSvalid, readingData, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      =      )           m_axis_tready : in  STD_LOGIC;�   	      =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   3   5          `                        m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   5   7          (                        bitCounter := 0;�   4   6          4                        state      <= waitingSvalid;5�_�   �   �           �   4   -    ����                                                                                                                                                                                                                                                                                                                            4   3       6   (       V   3    ^�     �   3   5   =      E                        m_axis_tvalid <= '0';--y ya no tengo mas nada5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            4   3       6   (       V   3    ^�     �   #   %   =    �   $   %   =    5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            5   3       7   (       V   3    ^�    �   #   %          +                        bitCounter    := 0;5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                               &          2       v   2    ^&    �         >      B   type shiftState is (waitingSvalid, readingData, waitingMready);5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                               &          2       v   2    ^�     �       "   >      !            s_axis_tready <= '0';5�_�   �   �           �   *        ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   *          F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);   y                        s_axis_tready              <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            *          *          V       ^�     �   (   +   <    �   )   *   <    5�_�   �   �           �   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �   +   ,          E                        bitCounter                 := bitCounter + 1;5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �   *   ,   =    �   +   ,   =    5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^�     �   )   *          y                        s_axis_tready              <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   +   #    ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^     �   *   ,   =      \                     if bitCounter < 8 then                             --porque bit voy?   5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^     �   +   ,                               else 5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^%     �   )   +          E                        bitCounter                 := bitCounter + 1;�   (   *          F                        m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^4     �   4   6   <    �   5   6   <    5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                            )   %       *   %       V   %    ^5     �   4   6          !            s_axis_tready <= '1';5�_�   �   �           �   4        ����                                                                                                                                                                                                                                                                                                                            4   *       4   *       V   *    ^:     �   3   4          7                        state         <= waitingSvalid;5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            4   *       4   *       V   *    ^:    �   5   7   <    �   6   7   <    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            4   *       4   *       V   *    ^     �   .   0   =    �   .   /   =    5�_�   �   �           �   .   $    ����                                                                                                                                                                                                                                                                                                                            5   *       5   *       V   *    ^"     �   .   0   >    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            6   *       6   *       V   *    ^#     �   /   1   ?    �   /   0   ?    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            7   *       7   *       V   *    ^$     �   .   0   @       5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            7   *       7   *       V   *    ^'     �   0   1          l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�   �   �           �   0   *    ����                                                                                                                                                                                                                                                                                                                            6   *       6   *       V   *    ^)     �   /   1   ?      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                            6   *       6   *       V   *    ^=    �       "   ?      !            s_axis_tready <= '1';5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /          0   %       V   %    ^�     �   .   /                               else   l                        s_axis_tready <= '1';                              --entonces yo tambien estoy listo5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                            /          /   %       V   %    ^�     �       "   =      !            s_axis_tready <= '0';5�_�   �   �           �   )   "    ����                                                                                                                                                                                                                                                                                                                            /          /   %       V   %    ^�     �   (   *   =      C                     m_axis_tdata(7-bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   )   "    ����                                                                                                                                                                                                                                                                                                                            /          /   %       V   %    ^�     �   (   *   =      B                     m_axis_tdata(-bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            )   ,       *   ,       V   ,    ^�    �   :   <   =         end process shift_reg;�   9   ;   =            end if;�   8   :   =               end if;�   7   9   =                  end case;�   6   8   =                        end if;�   5   7   =      7                        state         <= waitingSvalid;�   4   6   =      +                        bitCounter    := 0;�   3   5   =      -                        s_axis_tready <= '1';�   2   4   =      -                        m_axis_tvalid <= '0';�   1   3   =      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   0   2   =      $               when waitingMready =>�   /   1   =                        end if;�   .   0   =                           end if;�   -   /   =      7                        state         <= waitingMready;�   ,   .   =      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   +   -   =      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   *   ,   =      \                     if bitCounter = 8 then                             --porque bit voy?   �   )   +   =      @                     bitCounter               := bitCounter + 1;�   (   *   =      A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);�   '   )   =      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   =      $               when waitingSvalid =>�   %   '   =                  case state is�   $   &   =               else�   #   %   =                  bitCounter    := 0;�   "   $   =      -            m_axis_tdata  <= (others => '0');�   !   #   =      !            m_axis_tvalid <= '0';�       "   =      !            s_axis_tready <= '1';�      !   =      +            state         <= waitingSvalid;�          =               if rst = '0' then�         =            if rising_edge(clk) then�         =         begin�         =      0      variable bitCounter :integer range 0 to 8;�         =         shift_reg:process (clk) is�         =      ,   signal state:shiftState := waitingSvalid;�         =      5   type shiftState is (waitingSvalid, waitingMready);�         =      *           rst           : in  STD_LOGIC);�         =      )           clk           : in  STD_LOGIC;�         =      )           s_axis_tready : out STD_LOGIC;�         =      )           s_axis_tlast  : in  STD_LOGIC;�         =      )           s_axis_tvalid : in  STD_LOGIC;�         =      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      =      )           m_axis_tready : in  STD_LOGIC;�   	      =      )           m_axis_tlast  : out STD_LOGIC;�      
   =      )           m_axis_tvalid : out STD_LOGIC;�      	   =      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         =          Port(  �   (   *          A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);�   )   +          B                     bitCounter                 := bitCounter + 1;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^��    �                                      5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^��     �   (   +   =    �   )   *   =    5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            )          *                 ^��     �   '   )   ?      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            )          *                 ^��     �   )   +   ?      @                     bitCounter               := bitCounter + 1;�   (   *   ?      A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   +   #    ����                                                                                                                                                                                                                                                                                                                            )          *                 ^��     �   *   ,   ?    �   +   ,   ?    5�_�   �   �           �   ,   ,    ����                                                                                                                                                                                                                                                                                                                            )          *                 ^��     �   +   -   @      A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);5�_�   �   �           �   ,   ,    ����                                                                                                                                                                                                                                                                                                                            -   ?       -   ?       V   @    ^��     �   +   -   @      C                     m_axis_tdata(bitCounter_1) <= s_axis_tdata(0);5�_�   �   �           �   ,   @    ����                                                                                                                                                                                                                                                                                                                            -   ?       -   ?       V   @    ^��     �   +   -   @      C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(0);5�_�   �   �   �       �   +        ����                                                                                                                                                                                                                                                                                                                            ,   @       +   @       V   @    ^��     �   =   ?   @         end process shift_reg;�   <   >   @            end if;�   ;   =   @               end if;�   :   <   @                  end case;�   9   ;   @                        end if;�   8   :   @      7                        state         <= waitingSvalid;�   7   9   @      +                        bitCounter    := 0;�   6   8   @      -                        s_axis_tready <= '1';�   5   7   @      -                        m_axis_tvalid <= '0';�   4   6   @      �                  if m_axis_tready = '1' then                           --si el receptor puede recibir entonces ya latecho el dato..�   3   5   @      $               when waitingMready =>�   2   4   @                        end if;�   1   3   @                           end if;�   0   2   @      7                        state         <= waitingMready;�   /   1   @      `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   .   0   @      l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo�   -   /   @      \                     if bitCounter = 8 then                             --porque bit voy?   �   ,   .   @      @                     bitCounter               := bitCounter + 1;�   +   -   @      C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);�   *   ,   @      C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);�   )   +   @      B                     --bitCounter               := bitCounter + 1;�   (   *   @      C                     --m_axis_tdata(bitCounter) <= s_axis_tdata(0);�   '   )   @      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   @      $               when waitingSvalid =>�   %   '   @                  case state is�   $   &   @               else�   #   %   @                  bitCounter    := 0;�   "   $   @      -            m_axis_tdata  <= (others => '0');�   !   #   @      !            m_axis_tvalid <= '0';�       "   @      !            s_axis_tready <= '1';�      !   @      +            state         <= waitingSvalid;�          @               if rst = '0' then�         @            if rising_edge(clk) then�         @         begin�         @      0      variable bitCounter :integer range 0 to 8;�         @         shift_reg:process (clk) is�         @      ,   signal state:shiftState := waitingSvalid;�         @      5   type shiftState is (waitingSvalid, waitingMready);�         @      *           rst           : in  STD_LOGIC);�         @      )           clk           : in  STD_LOGIC;�         @      )           s_axis_tready : out STD_LOGIC;�         @      )           s_axis_tlast  : in  STD_LOGIC;�         @      )           s_axis_tvalid : in  STD_LOGIC;�         @      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   
      @      )           n_axis_tready : in  STD_LOGIC;�   	      @      )           m_axis_tlast  : out STD_LOGIC;�      
   @      )           m_axis_tvalid : out STD_LOGIC;�      	   @      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         @          Port(  �   *   ,          A                     m_axis_tdata(bitCounter) <= s_axis_tdata(0);�   +   -          C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);5�_�   �   �           �   +   >    ����                                                                                                                                                                                                                                                                                                                            ,   @       +   @       V   @    ^�      �   *   ,   @    �   +   ,   @    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            -   @       ,   @       V   @    ^�     �   *   ,   A      @                     bitCounter               := bitCounter + 1;5�_�   �   �           �   .   >    ����                                                                                                                                                                                                                                                                                                                            -   @       ,   @       V   @    ^�    �   -   /   A      @                     bitCounter               := bitCounter + 1;5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            )          +                 ^��     �   (   ,   A      C                     --m_axis_tdata(bitCounter) <= s_axis_tdata(0);   B                     --bitCounter               := bitCounter + 1;   B                     --bitCounter               := bitCounter + 1;5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            )          +                 ^��     �   *   +          @                     bitCounter               := bitCounter + 1;5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                            +          -          V       ^��    �   *   +          C                     m_axis_tdata(bitCounter)   <= s_axis_tdata(0);   C                     m_axis_tdata(bitCounter+1) <= s_axis_tdata(1);   @                     bitCounter               := bitCounter + 2;5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   
      =      )           n_axis_tready : in  STD_LOGIC;5�_�   �           �   �   +   @    ����                                                                                                                                                                                                                                                                                                                            ,   @       +   @       V   @    ^��     �   *   -   @      Aeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ceeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   -       ����                                                                                                                                                                                                                                                                                                                            0   *       0   *       V   *    ^A     �   ,   .   F      �                        state         <= readingData;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   q           s   r   (        ����                                                                                                                                                                                                                                                                                                                            0           1           V        ^ �     �   (   )   A    �   '   (   A      t                        m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   -           /   .      2    ����                                                                                                                                                                                                                                                                                                                               2          2       v   2    ^��     �         B      c--tomo 1 byte y mando 8 bytes en donde en cada unohhhhhhhhhhhhhhhhhhhhhhhhhhhde salida vale el bit05�_�   *           ,   +   *   &    ����                                                                                                                                                                                                                                                                                                                            <          <          V       ^�y     �   )   +   B      u                     state         <= ;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�                    2   G    ����                                                                                                                                                                                                                                                                                                                            1           2           V        ^�%     �   1   3   M      n                        bitCounter               := bitCounter+1;       hhhhhhhhhhhhhhhhhhhhhhhhhh--incremento5�_�                   1        ����                                                                                                                                                                                                                                                                                                                            1   #       2   #       V   #    ^�     �   0   3   M      Xeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�                    1   #    ����                                                                                                                                                                                                                                                                                                                            2   #       1   #       V   #    ^�     �   0   3   M      Xeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Teeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5��