Vim�UnDo� GwH�ddX
����ף�.��������ۙ��   )   entity lab1 is            �       �   �   �    ]���   H _�                            ����                                                                                                                                                                                                                                                                                                                                                             ]�>�     �               use IEEE.std_logic_1164.all.5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]�>�    �               use IEEE.std_logic_1164.all.;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]�>�    �                  N:=15�_�                    
   .    ����                                                                                                                                                                                                                                                                                                                                                             ]�>�    �   	            /      led: out std_logic_vector ( 3 downto 0 );5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�>�     �                  led(2)<=1;      led(3)<=0;�                  led(1)<=0;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�>�     �                  led(1)<=;0;      led(2)<=;1;      led(3)<=;0;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�>�    �                  led(2)<='1;      led(3)<='0;�                  led(1)<='0;5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             ]�s�     �                  led(0)<=swt(1);5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             ]�s�     �             �             5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             ]�s�     �             �             5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             ]�s�     �             �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�s�     �                  led(0)<=swt(0);�                  led(0)<=swt(0);�                  led(0)<=swt(0);�                  led(0)<=swt(0);5�_�                          ����                                                                                                                                                                                                                                                                                                                                                       ]�s�     �                  led(3)<=swt(0);�                  led(2)<=swt(0);�                  led(1)<=swt(0);�                  led(0)<=swt(0);5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]�s�    �                   led(1)<='0';      led(2)<='1';      led(3)<='0';5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�v+     �                  led(0)<=swt(0);      led(1)<=swt(1);      led(2)<=swt(2);      led(3)<=swt(3);5�_�                          ����                                                                                                                                                                                                                                                                                                                                                       ]�vN    �                  led(3)<=swt(3);�                  led(2)<=swt(3);�                  led(1)<=swt(3);�                  led(0)<=swt(3);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]��h     �                     �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]�È     �                  led(0)<=swt(3);      led(1)<=swt(2);      led(2)<=swt(1);      led(3)<=swt(0);5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]�Ì     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�â     �                        if(rst='1') then5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�ä     �                        if(rst='1'  then5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�æ     �                        elsif (clk=5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�ç     �                        elsif  clk=5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�ð     �                         elsif rising_edge( clk=5�_�                           ����                                                                                                                                                                                                                                                                                                                                                V       ]�ñ     �                        elsif rising_edge(clk=5�_�                       $    ����                                                                                                                                                                                                                                                                                                                                                V       ]�õ     �               %         elsif rising_edge(clk) then=5�_�                        #    ����                                                                                                                                                                                                                                                                                                                                                V       ]�ö     �                           �             5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                V       ]�ý     �                            if 5�_�       "           !           ����                                                                                                                                                                                                                                                                                                                                                V       ]�þ     �                   led(3)<=swt(0);�                   led(2)<=swt(1);�                   led(1)<=swt(2);�                   led(0)<=swt(3);5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �               /            led(0)<=            led(1)<=swt(2);�             �                           led(0)<=swt(3);               led(1)<=swt(2);5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �               5            led(0)<=led(3)            led(1)<=swt(2);5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �               6            led(0)<=led(3);            led(1)<=swt(2);5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �               ll            led(1)<=swt(2);5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �               l            led(1)<=swt(2);5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �             �             5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �             �             5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �             �             5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                v       ]���     �             �             5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                       ]���     �                           led(0)<=led(3);�                           led(0)<=led(3);�                           led(0)<=led(3);�                           led(0)<=led(3);5�_�   +   -           ,           ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                            led(0)<=led(3);               led(1)<=swt(2);               led(2)<=swt(1);               led(3)<=swt(0);5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                           led(1)<=led(3);5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                           led(2)<=led(3);5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                           led(3)<=led(3);5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                           led(3)<=led(1);5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                V       ]��
     �                           led(0)<=led(3);5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(1);5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(r);5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(r);5�_�   4   7           5          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(r);5�_�   5   8   6       7          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(r);5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led='0000'5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           �             5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                V       ]��<     �               	         �             5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                V       ]��B    �                        end if5�_�   ;   =           <   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]��d     �      
       �   	   
       5�_�   <   >           =   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]��e     �      
         /      swt: in  std_logic_vector ( 3 downto 0 );5�_�   =   ?           >   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �      
         /      clk: in  std_logic_vector ( 3 downto 0 );5�_�   >   @           ?   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �      
         '      clk: in  std_logic( 3 downto 0 );5�_�   ?   A           @   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �      
       �   	   
       5�_�   @   B           A   	       ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �      
               clk: in  std_logic;5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                V       ]���   	 �                	         �             5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                         if rst='1'  then5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                V       ]���   
 �                            led='0001'5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �                            led<='0001'5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                                V       ]��:    �                            led<='0001';5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                V       ]��E     �                            led<='0001'5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                V       ]��F    �                            led<="0001'5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                V       ]��G    �                            led<="0001"5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                                                V       ]��O    �                            led<="0001";5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                V       ]��Z    �                            led<="0001"5�_�   K   N           L          ����                                                                                                                                                                                                                                                                                                                                                V       ]�ƛ     �              5�_�   L   O   M       N          ����                                                                                                                                                                                                                                                                                                                                                  V       ]�ơ     �         "      	         �         !    5�_�   N   P           O      	    ����                                                                                                                                                                                                                                                                                                                            !          !          V       ]���     �         "               variable i:=05�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                            !          !          V       ]���     �         "      "         signal led0;variable i:=05�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                                       ]���     �         "                  led(1)<=led(2);               led(2)<=led(3);               led(3)<=led(0);�         "                  led(0)<=led(1);5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                                       ]���    �         "                  led(0)<='1'led(1);               led(1)<='1'led(2);               led(2)<='1'led(3);               led(3)<='1'led(0);5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �                         signal led0;5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �         !    �         !    5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �         "               signal led0;5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �         "      ,         signal led0: std_logic(0 downto 0);5�_�   V   X           W           ����                                                                                                                                                                                                                                                                                                                                                             ]�F�     �         "         begin5�_�   W   Y           X           ����                                                                                                                                                                                                                                                                                                                                                             ]�F�     �                 5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(1)<='1';               led(2)<='1';               led(3)<='1';�         !                  led(0)<='1';5�_�   Y   ^           Z          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(0)<=led(3)'1';               led(1)<=led(3)'1';               led(2)<=led(3)'1';               led(3)<=led(3)'1';5�_�   Z   _   [       ^          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(0)<=led(3)';               led(1)<=led(3)';               led(2)<=led(3)';               led(3)<=led(3)';5�_�   ^   a           _          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�    �         !                  led(3)<=led(3);�         !                  led(2)<=led(3);�         !                  led(1)<=led(3);�         !                  led(0)<=led(3);5�_�   _   b   `       a          ����                                                                                                                                                                                                                                                                                                                                                             ]�Gk     �         !      ,         signal led0: std_logic(3 downto 0);5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                                             ]�Gm     �         !      /         signal led_in0: std_logic(3 downto 0);5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                                       ]�Gu     �         !                  led(1)<=led(2);               led(2)<=led(1);               led(3)<=led(0);�         !                  led(0)<=led(3);5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                       ]�G�     �         "                  �         !    5�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                                                       ]�G�     �                            led_in5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                                                       ]�G�    �         !       5�_�   f   i           g      !    ����                                                                                                                                                                                                                                                                                                                                                       ]�G�    �         !      .         signal led_in: std_logic(3 downto 0);5�_�   g   j   h       i          ����                                                                                                                                                                                                                                                                                                                            	           
           V        ]�I�     �         !    �         !    5�_�   i   l           j          ����                                                                                                                                                                                                                                                                                                                            	           
           V        ]�I�    �         "                  led<="0001";5�_�   j   m   k       l           ����                                                                                                                                                                                                                                                                                                                                                V       ]�I�     �      !   "            end process;�          "               end if;�         "                  led(3)<=led_in(0);�         "                  led(2)<=led_in(1);�         "                  led(1)<=led_in(2);�         "                  led(0)<=led_in(3);�         "      $         elsif rising_edge(clk) then�         "                  led_in <= "0001";�         "                  led    <= "0001";�         "               if rst<='1'  then�         "            begin�         "            process(clk,rst)�         "         begin�         "      5         signal led_in: std_logic_vector(3 downto 0);�         "          );�         "      .      led: out std_logic_vector ( 3 downto 0 )�   
      "      /      swt: in  std_logic_vector ( 3 downto 0 );�   	      "            clk: in  std_logic;�      
   "            rst: in  std_logic;�      	   "      	   port (�         "         );�         "         N: natural :=1�         "         generic (�                            led<="0001";�                            led_in<="0001";5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                                V       ]�I�     �         "                  led    <= "0001";5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                                                V       ]�I�     �          #                  �          "    5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                                                       ]�I�     �         #                  led(1)<=led_in(2);               led(2)<=led_in(1);               led(3)<=led_in(0);�         #                  led(0)<=led_in(3);5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                                                       ]�I�    �          #                  led<=led_in5�_�   p   r           q          ����                                                                                                                                                                                                                                                                                                                                                       ]�K�     �         #               if rst<='1'  then5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                                                       ]�K�    �         #               if rst=='1'  then5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                                                       ]�K�    �         #               if rst='1'  then5�_�   s   u           t          ����                                                                                                                                                                                                                                                                                                                                                       ]�L~     �         #      !            led_in(0)<=led_in(3);   !            led_in(1)<=led_in(2);   !            led_in(2)<=led_in(1);   !            led_in(3)<=led_in(0);5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                       ]�L�     �         #      !            led_in(3)<=led_in(1);�         #      !            led_in(2)<=led_in(1);�         #      !            led_in(1)<=led_in(1);�         #      !            led_in(0)<=led_in(1);5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                                                       ]�L�    �         #      !            led_in(3)<=led_in(4);5�_�   v   x           w           ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�L�     �                            led<=led_in;5�_�   w   y           x       	    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�L�     �      !   "    �       !   "    5�_�   x   z           y           ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�L�     �      !                      led<=led_in;5�_�   y   {           z            ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M     �                          led<=led_in;5�_�   z   |           {   !       ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M   ! �       "   "    �   !   "   "    5�_�   {   }           |   !   	    ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M   " �       "                   led<=led_in;5�_�   |   ~           }           ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M4   # �                 5�_�   }              ~      	    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�Mb     �                5         signal led_in: std_logic_vector(3 downto 0);5�_�   ~   �                 .    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�M�   $ �         "      /   signal led_in: std_logic_vector(3 downto 0);5�_�      �           �      /    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�M�     �         "      6   signal led_in: std_logic_vector(3 downto 0)='0000';5�_�   �   �   �       �      4    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�N   % �         "      6   signal led_in: std_logic_vector(3 downto 0)="0000';5�_�   �   �           �      .    ����                                                                                                                                                                                                                                                                                                                               	          	       V   	    ]�N   & �         "      6   signal led_in: std_logic_vector(3 downto 0)="0000";5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                                                  V       ]�N     �                       led<=led_in;5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                                                  V       ]�N#     �      !   !    �       !   !    5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                                                  V       ]�N'     �                       led<=led_in;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V       ]�N)   ( �          !    �          !    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�N}     �                      led<=led_in;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�N   ) �      !   !    �       !   !    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�N�   * �         "                  led    <= "0000";5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�N�   + �                      --      led    <= "0000";5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�Tn   , �   
      !      /      swt: in  std_logic_vector ( 3 downto 0 );5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�XW     �   
      !      1--      swt: in  std_logic_vector ( 3 downto 0 );5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�XW     �   
      !      0-      swt: in  std_logic_vector ( 3 downto 0 );5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                V       ]�XX   - �   
      !      /      swt: in  std_logic_vector ( 3 downto 0 );5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�X`     �         !            process(clk,rst)5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�Xl     �         !      $         elsif rising_edge(clk) then5�_�   �   �           �      !    ����                                                                                                                                                                                                                                                                                                                                                V       ]�Xs   . �         !      *         elsif rising_edge(swt(0)clk) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�[     �         !            process(clk,swt(0))5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�[    0 �         !            process(swt(0))5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                             ]�dQ     �         !      '         elsif rising_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ]�dT     �         !    �         !    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ]�dU     �         "      )--         elsif rising_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ]�dV     �         "      (-         elsif rising_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ]�dY     �         "      '         elsif rising_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ]�dY   1 �         "               els5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ]�e-     �         "               else5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             ]�e-     �         "               els5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                             ]�e.     �                         el5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ]�e1     �         !      )--         elsif rising_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             ]�e1     �         !      (-         elsif rising_edge(swt(0)) then5�_�   �   �           �      !    ����                                                                                                                                                                                                                                                                                                                                                v       ]�ep     �         !      '         elsif rising_edge(swt(0)) then5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�ey     �         !      '         elsif rising_edge(swt(0)) then5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�e|     �         !      +         elsif rising_edge(swt(0)) or  then�         !    5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�e~   2 �         !      >         elsif rising_edge(swt(0)) or rising_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�f�   3 �         !      ?         elsif rising_edge(swt(0)) or falling_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�f�     �         "                  �         !    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�f�   4 �         "               end if;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�g^     �         "      A--         elsif rising_edge(swt(0)) or falling_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�g^     �         "      @-         elsif rising_edge(swt(0)) or falling_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�ga     �         "      ?         elsif rising_edge(swt(0)) or falling_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�gc     �         "      ?         elsif rising_edge(clk(0)) or falling_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�gc     �         "      >         elsif rising_edge(clk0)) or falling_edge(swt(0)) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         !       v   !    ]�gc     �         "      =         elsif rising_edge(clk)) or falling_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                          6       v   6    ]�gh     �         "      <         elsif rising_edge(clk) or falling_edge(swt(0)) then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                          6       v   6    ]�gi     �         "      %         elsif rising_edge(clk)  then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                          6       v   6    ]�gk     �         #                  �         "    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                          6       v   6    ]�gz     �          $                  �          #    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         $            process(rst,swt(0))5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         $            process(rst,clk))5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �                         end if;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         $         �         #    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         %                     �         $    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �      "   &                  �      !   %    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                  if(swt(0)=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                  if (swt(0)=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                  if swt(0)=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                     latch:=15�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                     latch:=1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                    latch:=1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]�g�     �         '                   latch:=1;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�g�     �      !                   else�                 !            led_in(3)<=led_in(0);�                !            led_in(2)<=led_in(3);�                !            led_in(1)<=led_in(2);�                !            led_in(0)<=led_in(1);�                            latch:=1;5�_�   �   �           �   "   	    ����                                                                                                                                                                                                                                                                                                                                                 V       ]�g�     �   !   "                   else5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                                 V       ]�g�     �   !   #   &      --         end if;5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                                 V       ]�g�     �   !   #   &      -         end if;5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                            "                     V       ]�g�     �   !   #                   end if;�       "                      latch=0;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                      #          V       ]�g�   5 �   "   $                end process;5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                      #          V       ]�g�     �   "   $   &               end process;5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                      #          V       ]�g�     �   "   $   &              end process;5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                      #          V       ]�g�   7 �   "   $   &             end process;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�h     �                    variable latch: unsigned :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�h   8 �         %    �         %    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�h     �                    variable latch: unsigned :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�h     �         %    �         %    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�h    9 �                    variable latch: unsigned :=0;5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                                V       ]�h+   : �       "   &                     latch=0;5�_�   �   �           �   "   
    ����                                                                                                                                                                                                                                                                                                                                                V       ]�h4   ; �   "   $   '                  �   "   $   &    5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                                V       ]�h9   = �   "   $   '               end if;;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�h�   > �         '      &         variable latch: unsigned :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�h�     �         '      )            if swt(0)=0  and latch=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�h�     �         '      )            if swt(0)=0  and latch=0 then5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�h�     �         '      *            if swt(0)='0  and latch=0 then5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�h�   @ �         '      *            if swt(0)='0' and latch=0 then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�iW     �         '      %         variable latch: integer :=0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�iX     �         '      $         variable latch: integer:=0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�iX     �         '      #         variable latch: integer=0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $                    V       ]�iX   A �         '      "         variable latch: integer0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i{     �         '      *            if swt(0)='0' and latch=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i|     �         (                     �         '    5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i�     �         (                     if 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i�     �                               latch:=1;5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �      !          $               led_in(3)<=led_in(0);�                 $               led_in(2)<=led_in(3);�                $               led_in(1)<=led_in(2);�                $               led_in(0)<=led_in(1);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �       "   )                        �       "   (    5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   !   "                      else5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   !   #                         latch:=0;5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �       "   )                        �       "   (    5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   !   #                         else5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   "   $                            latch:=0;5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�   B �   #   $                      end if;5�_�   �   �   �       �   $       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   #   %   (    �   $   %   (    5�_�   �   �   �       �   $        ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]�i�   C �   #   %                   end if;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )                     if latch=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )                     if latch>=0 then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )                        latch:=1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )      $                  latch:=latcj-1hh1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )      $                  latch:=latch-1hh1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��     �         )      #                  latch:=latch-hh1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��      �         )      "                  latch:=latch-h1;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]��!     �         *                        �         )    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            '   	          	       V   	    ]��.     �         *    �         *    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ]��2     �         +      !                  latch:=latch-1;5�_�   �   �           �   $        ����                                                                                                                                                                                                                                                                                                                            $          %          V       ]��A   D �   #   $                      else                  latch:=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]���     �         )      !                  latch:=5000000;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]���   G �         )      $                  latch:=1005000000;5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]���   H �         )      entity lab1 is5�_�   �           �   �           ����                                                                                                                                                                                                                                                                                                                            &   	          	       V   	    ]�i�     �                '            if swt(0)        = '0' then�                %               if latch      = 0 then�                !                  latch     := 1;�                )                  led_in(0) <= led_in(1);�   "   $          !               latch        := 0;�      !          )                  led_in(3) <= led_in(0);�                 )                  led_in(2) <= led_in(3);�                (         if rst              = '1'  then�                &            led_in          <= "0001";�                )                  led_in(1) <= led_in(2);�         )         generic (�         )         N: natural :=1�         )         );�      	   )      	   port (�      
   )            rst: in  std_logic;�   	      )            clk: in  std_logic;�   
      )      /      swt: in  std_logic_vector ( 2 downto 0 );�         )      .      led: out std_logic_vector ( 3 downto 0 )�         )          );�         )      7   signal led_in: std_logic_vector(3 downto 0):="0000";�         )         begin�         )            process(rst,clk)�         )      !         variable latch: integer;�         )            begin�         )      (         if rst              = '1'  then�         )      &            led_in          <= "0001";�         )      $         elsif rising_edge(clk) then�         )      '            if swt(0)        = '0' then�         )      %               if latch      = 0 then�         )      !                  latch     := 1;�         )      )                  led_in(0) <= led_in(1);�         )      )                  led_in(1) <= led_in(2);�          )      )                  led_in(2) <= led_in(3);�      !   )      )                  led_in(3) <= led_in(0);�       "   )                     end if;�   !   #   )                  else�   "   $   )      !               latch        := 0;�   #   %   )               end if;�   $   &   )               end if;�   %   '   )            end process;�   &   (   )            led<=led_in;5�_�   �           �   �   "       ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �   "   #   (       5�_�   �           �   �           ����                                                                                                                                                                                                                                                                                                                                                 V       ]�i�     �       !   (    �       !   (                  else5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i�     �         (    �         (      '                  land latch=0 atch:=1;5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                         %       v   %    ]�i�     �         (                     if latch:=1;5�_�   �       �   �   �          ����                                                                                                                                                                                                                                                                                                                            %                    V       ]�h�     �         '                  if swt(0)='0               and latch=0 then5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                            %                    V       ]�h�     �         '                  if swt(0)='0               and latch=0 then5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                                             ]�dG     �         !      &         else rising_edge(swt(0)) then5�_�   �       �   �   �      0    ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M�     �         "      0   signal led_in: std_logic_vector(3 downto 0)="      000';5�_�   �           �   �      0    ����                                                                                                                                                                                                                                                                                                                                	           	       V   	    ]�M�     �         "      0   signal led_in: std_logic_vector(3 downto 0)="      000';5�_�   j           l   k           ����                                                                                                                                                                                                                                                                                                                                                V       ]�I�     �         "      eeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   g           i   h      4    ����                                                                                                                                                                                                                                                                                                                            	           
           V        ]�I�     �         !      7         signal led_in: std_logic_vector(3 downto 0):=;5�_�   _           a   `      .    ����                                                                                                                                                                                                                                                                                                                                                             ]�G     �   
      !      .      swt: in  std_logic_vector ( 3 downto 0 )5�_�   Z   \       ^   [          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(3)<=led(3);5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(0)<=led(3)';�         !                  led(1)<=led(3)';�         !                  led(2)<=led(3)';�         !                  led(3)<=led(3);5�_�   \               ]          ����                                                                                                                                                                                                                                                                                                                                                       ]�F�     �         !                  led(0)<=led(3)';�         !                  led(1)<=led(4)';�         !                  led(2)<=led(5)';�         !                  led(3)<=led(6);5�_�   L           N   M          ����                                                                                                                                                                                                                                                                                                                                                  V       ]�ƞ     �         !    �         !            process;(clk,rst)5�_�   5           7   6          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                           led(2)<=led(3335�_�                          ����                                                                                                                                                                                                                                                                                                                                                       ]�vF     �                  led(0)<=swt(3);�                  led(1)<=swt(4);�                  led(2)<=swt(5);�                  led(3)<=swt(6);5�_�                          ����                                                                                                                                                                                                                                                                                                                                                       ]�v?     �                  led(0)<=swt(3);�                  led(1)<=swt(4);�                  led(2)<=swt(5);�                  led(3)<=swt(6);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�v3     �                  led(0)<=swt(3);�                  led(1)<=swt(4);�                  led(2)<=swt(5);�                  led(3)<=swt(6);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ]�s�     �             �                  led(0)<=swt(0);5��