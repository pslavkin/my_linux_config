Vim�UnDo� ����4�t*f���hq�Ґ�c����%���   A                                   ^O    _�                              ����                                                                                                                                                                                                                                                                                                                                                             ^N    �                (architecture Behavioral of split_2to8 is�                end split_2to8;�                entity split_2to8 is5��