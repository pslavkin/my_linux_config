Vim�UnDo� ��/� K��������Q%oX1Y94��㎤   ?   C                        m_axis_tdata  <= s_axis_tdata(15 downto 8);   3   6      #       #   #   #    ^d�    _�                             ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �                *architecture Behavioral of slice_2from8 is�                end slice_2from8;�                entity slice_2from8 is5�_�                    +   !    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   *   ,   A      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    +   !    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   *   ,   A      S                     m_axis_tdata0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    +   !    ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �   *   ,   A      R                     m_axis_tdata) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    +   2    ����                                                                                                                                                                                                                                                                                                                                                v       ^�#     �   *   ,   A      Q                     m_axis_tdata <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    +   >    ����                                                                                                                                                                                                                                                                                                                                                v       ^�D     �   *   ,   A      Q                     m_axis_tdata <= s_axis_tdata(7 downto 0);    --pongo el dato5�_�      	              ,       ����                                                                                                                                                                                                                                                                                                                                                v       ^�E     �   +   ,          V                     m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�      
          	   )        ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�O     �   =   ?   @         end process shift_reg;�   <   >   @            end if;�   ;   =   @               end if;�   :   <   @                  end case;�   9   ;   @                        end if;�   8   :   @                           end if;�   7   9   @      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   6   8   @      -                        s_axis_tready <= '1';�   5   7   @      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   4   6   @                           else�   3   5   @      Y                        m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato�   2   4   @      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato�   1   3   @      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   0   2   @      Q                     bitCounter := bitCounter+2;                     --incremento�   /   1   @      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?�   .   0   @      $               when waitingMready =>�   -   /   @                        end if;�   ,   .   @      }                     state         <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   +   -   @      o                     m_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   *   ,   @      ?                     m_axis_tdata  <= s_axis_tdata(7 downto 0);�   )   +   @      (                     bitCounter    := 0;�   (   *   @      *                     s_axis_tready <= '0';�   '   )   @      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   &   (   @      $               when waitingSvalid =>�   %   '   @                  case state is�   $   &   @               else�   #   %   @      -            m_axis_tdata  <= (others => '0');�   "   $   @      !            m_axis_tvalid <= '0';�   !   #   @      !            s_axis_tready <= '1';�       "   @      +            state         <= waitingSvalid;�      !   @               if rst = '0' then�          @            if rising_edge(clk) then�         @         begin�         @      0      variable bitCounter :integer range 0 to 8;�         @         shift_reg:process (clk) is�         @      ,   signal state:shiftState := waitingSvalid;�         @      5   type shiftState is (waitingSvalid, waitingMready);�         @      *           rst           : in  STD_LOGIC);�         @      )           clk           : in  STD_LOGIC;�         @      )           s_axis_tready : out STD_LOGIC;�         @      )           s_axis_tlast  : in  STD_LOGIC;�         @      )           s_axis_tvalid : in  STD_LOGIC;�         @      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         @      )           m_axis_tready : in  STD_LOGIC;�   
      @      )           m_axis_tlast  : out STD_LOGIC;�   	      @      )           m_axis_tvalid : out STD_LOGIC;�      
   @      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      	   @          Port(  �   (   *          ,                     s_axis_tready   <= '0';�   ,   .                               state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   +   -          q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato�   *   ,          >                     m_axis_tdata <= s_axis_tdata(7 downto 0);�   )   +          *                     bitCounter      := 0;5�_�   	              
   1   .    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�[     �   0   2   @      Q                     bitCounter := bitCounter+2;                     --incremento5�_�   
                 2   #    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�^     �   1   3   @      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�                    3   #    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�m     �   2   4   @    �   3   4   @    5�_�                    3       ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�o     �   2   4          ?                     m_axis_tdata  <= s_axis_tdata(7 downto 0);5�_�                    2   %    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�p     �   1   3   A      f                     if bitCounter = 8 then                             --perfecto, porque bit voy?   5�_�                    3   6    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�v     �   2   4   A      B                        m_axis_tdata  <= s_axis_tdata(7 downto 0);5�_�                    3   @    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�z     �   2   4   A      C                        m_axis_tdata  <= s_axis_tdata(15 downto 0);5�_�                    3   @    ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�z     �   2   4   A      C                        m_axis_tdata  <= s_axis_tdata(15 downto 9);5�_�                    4        ����                                                                                                                                                                                                                                                                                                                            4   ?       5   ?       V   ?    ^�|    �   3   4          W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato   Y                        m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�                   	   1    ����                                                                                                                                                                                                                                                                                                                                                             ^�7     �      
   ?      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�                       1    ����                                                                                                                                                                                                                                                                                                                                                             ^�@    �         ?      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�                       1    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �         ?      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);5�_�                       .    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �         ?      0      variable bitCounter :integer range 0 to 8;5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �         ?      2      variable bitCounter :integer range 0 to 488;5�_�                    1   .    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   0   2   ?      Q                     bitCounter := bitCounter+1;                     --incremento5�_�                    2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter = 1 then                             --perfecto, porque bit voy?   5�_�                    2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter m 1 then                             --perfecto, porque bit voy?   5�_�                    2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter , 1 then                             --perfecto, porque bit voy?   5�_�                    2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter m 1 then                             --perfecto, porque bit voy?   5�_�                    2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter m 1 then                             --perfecto, porque bit voy?   5�_�                     2   #    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter M 1 then                             --perfecto, porque bit voy?   5�_�      !               2   %    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   1   3   ?      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   5�_�       "           !   3   6    ����                                                                                                                                                                                                                                                                                                                                                             ^c�     �   2   4   ?      C                        m_axis_tdata  <= s_axis_tdata(15 downto 8);5�_�   !   #           "   3   J    ����                                                                                                                                                                                                                                                                                                                                                             ^c�    �   2   4   ?      M                        m_axis_tdata  <= s_axis_tdata(bitCounter+8 downto 8);5�_�   "               #   3   A    ����                                                                                                                                                                                                                                                                                                                                                             ^d�    �   2   4   ?      V                        m_axis_tdata  <= s_axis_tdata(bitCounter+8 downto bitCounter);5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            4   ?       4   ?       V   ?    ^�~     �   3   5        5�_�              	      )        ����                                                                                                                                                                                                                                                                                                                            )          -          V       ^�M     �   (   .   @      ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   >eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   qeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5��