Vim�UnDo� f�K:����!�xU���	 �9L'7u�sg���7W   )   :           inData   : in    std_logic_vector (7 downto 0),   
   9      �   �   �   �   �    ]���   + _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ]��m     �                 R----------------------------------------------------------------------------------   -- Company:    -- Engineer:    --    &-- Create Date: 12/04/2019 04:59:29 PM   -- Design Name:    #-- Module Name: spi28b - Behavioral   -- Project Name:    -- Target Devices:    -- Tool Versions:    -- Description:    --    -- Dependencies:    --    -- Revision:   -- Revision 0.01 - File Created   -- Additional Comments:   --    R----------------------------------------------------------------------------------        5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  V        ]��p     �                    7-- Uncomment the following library declaration if using   6-- arithmetic functions with Signed or Unsigned values5�_�                            ����                                                                                                                                                                                                                                                                                                                                       	           V        ]��|    �                ?-- Uncomment the following library declaration if instantiating   &-- any Xilinx leaf cells in this code.   --library UNISIM;   --use UNISIM.VComponents.all;    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]���     �         2      D    signal bitCount   : std_logic_vector (7 downto 0) := "00000001";5�_�                           ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]���     �         2      6    signal bitCount   : in (7 downto 0) := "00000001";5�_�                           ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]���     �         2      8    variable bitCount   : in (7 downto 0) := "00000001";5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]���     �         2      A    variable bitCount   : integer lin (7 downto 0) := "00000001";5�_�      	                 )    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]���     �         2      C    variable bitCount   : integer range (7 downto 0) := "00000001";5�_�      
           	      )    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      C    variable bitCount   : integer range (8 downto 0) := "00000001";5�_�   	              
      )    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      C    variable bitCount   : integer range (9 downto 0) := "00000001";5�_�   
                    +    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      C    variable bitCount   : integer range (0 downto 0) := "00000001";5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      B    variable bitCount   : integer range (0 ownto 0) := "00000001";5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      A    variable bitCount   : integer range (0 wnto 0) := "00000001";5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      @    variable bitCount   : integer range (0 nto 0) := "00000001";5�_�                       .    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      ?    variable bitCount   : integer range (0 to 0) := "00000001";5�_�                       (    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      ?    variable bitCount   : integer range (0 to 8) := "00000001";5�_�                       .    ����                                                                                                                                                                                                                                                                                                                                         	       v   	    ]��     �         2      >    variable bitCount   : integer range 0 to 8) := "00000001";5�_�                       2    ����                                                                                                                                                                                                                                                                                                                               2          ;       v   ;    ]��     �         2      =    variable bitCount   : integer range 0 to 8 := "00000001";5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            "          "   '       v   '    ]��     �   !   #   2      A                    bitCount(7 downto 1) <= bitCount(6 downto 0);5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            "          "   '       v   '    ]��     �   !   #   2      5                    bitCount <= bitCount(6 downto 0);5�_�                    "       ����                                                                                                                                                                                                                                                                                                                            "          "   '       v   '    ]��     �   !   #   2      6                    bitCount :<= bitCount(6 downto 0);5�_�                    "   (    ����                                                                                                                                                                                                                                                                                                                            "   (       "   3       v   3    ]��     �   !   #   2      5                    bitCount := bitCount(6 downto 0);5�_�                    $   #    ����                                                                                                                                                                                                                                                                                                                            $   #       $   ,       v   ,    ]��&    �   #   %   2      3                    if (bitCount = "00000000") then5�_�                    )   %    ����                                                                                                                                                                                                                                                                                                                            )   %       )   .       v   .    ]��:    �   (   *   2      0                        bitCount   <="00000001";5�_�                           ����                                                                                                                                                                                                                                                                                                                            )   %       )   .       v   .    ]��K     �         2      4    variable bitCount   : integer range 0 to 8 := 0;5�_�                           ����                                                                                                                                                                                                                                                                                                                            )   %       )   .       v   .    ]��K     �         2      3    variable bitCount  : integer range 0 to 8 := 0;5�_�                       '    ����                                                                                                                                                                                                                                                                                                                            )   %       )   .       v   .    ]��N    �         2      2    variable bitCount : integer range 0 to 8 := 0;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]��Y     �                2    variable bitCount : integer range 0 to 8 := 0;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]��^     �         1    �         1    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                V       ]��`    �                 5�_�                     (   #    ����                                                                                                                                                                                                                                                                                                                                                V       ]��k    �   '   )   1      (                        bitCount   <= 0;5�_�      !               ,       ����                                                                                                                                                                                                                                                                                                                                                V       ]��q     �   +   -   1      *                  bitCount   <="00000001";5�_�       "           !   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]��s     �   +   -   1      *                  bitCount   :="00000001";5�_�   !   #           "   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]��t     �   +   -   1      #                  bitCount   :=01";5�_�   "   $           #   ,   !    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]��u     �   +   -   1      $                  bitCount   := 01";5�_�   #   %           $   ,   !    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]��u    �   +   -   1      #                  bitCount   := 0";5�_�   $   &           %   0        ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�K     �   /   1   1       5�_�   %   '           &   0       ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�Y     �   /   0             bitCount_sig <= bitCount;5�_�   &   (           '   (   #    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�^     �   '   )   0      (                        bitCount   := 0;5�_�   '   )           (   (   &    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�b     �   '   )   0      (                        bitCount   <= 0;5�_�   (   *           )   (   (    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�d     �   '   )   0      )                        bitCount   <= "0;5�_�   )   +           *   #   #    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�m     �   "   $   0      *                    if (bitCount = 8) then5�_�   *   ,           +   #   (    ����                                                                                                                                                                                                                                                                                                                            ,          ,   %       v   %    ]�t     �   "   $   0      /                    if (bitCount = "100"8) then5�_�   +   -           ,   (   '    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]�v     �   '   )   0      1                        bitCount   <= "00000000";5�_�   ,   .           -   #   $    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]�|     �   "   $   0      .                    if (bitCount = "100") then5�_�   -   /           .   #   &    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]�~     �   "   $   0      0                    if (bitCount = "10100") then5�_�   .   0           /   !       ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]��     �       "   0      -                    bitCount := bitCount + 1;5�_�   /   1           0   !        ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]��     �       "   0      -                    bitCount <= bitCount + 1;5�_�   0   2           1   !   1    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]��     �       "   0      >                    bitCount <= std_logic_vector(bitCount + 1;5�_�   1   3           2   !   B    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]��     �       "   0      G                    bitCount <= std_logic_vector(unsigned(bitCount + 1;5�_�   2   4           3   !   G    ����                                                                                                                                                                                                                                                                                                                            (   '       (   +       v   +    ]��     �       "   0      H                    bitCount <= std_logic_vector(unsigned(bitCount) + 1;5�_�   3   5           4           ����                                                                                                                                                                                                                                                                                                                               1          1       V   G    ]��     �                2    variable bitCount : integer range 0 to 8 := 0;5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                               1          1       V   G    ]��     �         /    �         /    5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                               1          1       V   G    ]��     �         0      2    variable bitCount : integer range 0 to 8 := 0;5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                               1          1       V   G    ]��     �         0      1    signal  bitCount : integer range 0 to 8 := 0;5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                               1          1       V   G    ]��     �         0      0    signal bitCount : integer range 0 to 8 := 0;5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                v       ]��     �         0      2    signal bitCount   : integer range 0 to 8 := 0;�         0    5�_�   9   ;           :      )    ����                                                                                                                                                                                                                                                                                                                                         '       v       ]��     �         0      ;    signal bitCount   : std_logic_vector range 0 to 8 := 0;5�_�   :   <           ;      I    ����                                                                                                                                                                                                                                                                                                                                         '       v       ]��    �         0      [    signal bitCount   : std_logic_vector (3 downto 0) := (others => '0');range 0 to 8 := 0;5�_�   ;   =           <           ����                                                                                                                                                                                                                                                                                                                                                V   H    ]��     �                                                          5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                V   H    ]��     �                                    5�_�   =   @           >          ����                                                                                                                                                                                                                                                                                                                                                V   H    ]��     �                                    5�_�   >   A   ?       @           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   *   ,   ,              end process;�   )   +   ,                   end if;�   (   *   ,                      end if;�   '   )   ,      "                  bitCount   := 0;�   &   (   ,                      else �   %   '   ,                          end if;�   $   &   ,                              �   #   %   ,      ,                        bitCount   <= "000";�   "   $   ,      =                        ledsData   <= mosiSignal(3 downto 0);�   !   #   ,      1                        outData    <= mosiSignal;�       "   ,      4                        spi_miso   <= misoSignal(7);�      !   ,      -                        misoSignal <= inData;�          ,      /                    if (bitCount = "1000") then�         ,      W                    bitCount               <= std_logic_vector(unsigned(bitCount) + 1);�         ,      E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);�         ,      <                    spi_miso               <= misoSignal(7);�         ,      7                    mosiSignal(0)          <= spi_mosi;�         ,      E                    mosiSignal(7 downto 1) <= mosiSignal(6 downto 0);�         ,      "                if (cs = '0') then�         ,      $            if rising_edge(clk) then�         ,              begin�         ,          process (clk)�         ,      begin   �         ,      I    signal bitCount   : std_logic_vector (3 downto 0) := (others => '0');�         ,      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         ,      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         ,      '           clk      : in    STD_LOGIC);�   
      ,      :           ledsData : out   std_logic_vector (3 downto 0);�   	      ,      :           inData   : in    std_logic_vector (7 downto 0);�      
   ,      :           outData  : out   std_logic_vector (7 downto 0);�      	   ,      &           cs       : in    std_logic;�         ,      &           spi_miso : out   STD_LOGIC;�         ,      &    Port ( spi_mosi : in    STD_LOGIC;�                E                    mosiSignal(7 downto 1) <= mosiSignal(6 downto 0);�                I                    bitCount <= std_logic_vector(unsigned(bitCount) + 1);�                E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);�                .                    spi_miso <= misoSignal(7);�                .                    mosiSignal(0) <= spi_mosi;5�_�   @   B           A   $   '    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   #   %   ,      ,                        bitCount   <= "000";5�_�   A   C           B   (       ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   '   )   ,      "                  bitCount   := 0;5�_�   B   D           C   (       ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   '   )   ,      #                  bitCount   <:= 0;5�_�   C   E           D   (        ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   '   )   ,      "                  bitCount   <= 0;5�_�   D   F           E   (   %    ����                                                                                                                                                                                                                                                                                                                                                V       ]��   	 �   '   )   ,      &                  bitCount   <= "0000;5�_�   E   G           F      $    ����                                                                                                                                                                                                                                                                                                                                                V       ]�0     �          ,      /                    if (bitCount = "1000") then5�_�   F   H           G      %    ����                                                                                                                                                                                                                                                                                                                                                V       ]�1   
 �          ,      /                    if (bitCount = "0000") then5�_�   G   I           H      $    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �          ,      /                    if (bitCount = "0111") then5�_�   H   J           I   $   '    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   #   %   ,      -                        bitCount   <= "0000";5�_�   I   K           J      *    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         ,      I    signal bitCount   : std_logic_vector (3 downto 0) := (others => '0');5�_�   J   L           K   (   #    ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �   '   )   ,      '                  bitCount   <= "0000";5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �         ,    5�_�   L   N           M      D    ����                                                                                                                                                                                                                                                                                                                                                V       ]�Y     �         -      E                    mosiSignal(7 downto 1) <= mosiSignal(6 downto 0);5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]�e     �         -      P                    mosiSignal(7 downto 1) <= mosiSignal(6 downto 0) & spi_mosi;5�_�   N   P           O          ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]�h    �         -      7                    mosiSignal(0)          <= spi_mosi;5�_�   O   Q           P      -    ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]�t     �         -      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   P   R           Q      6    ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]�v     �         -      D                    mosiSignal <= mosiSignal(7 downto 0) & spi_mosi;5�_�   Q   S           R      -    ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��     �         -      D                    mosiSignal <= mosiSignal(7 downto 1) & spi_mosi;5�_�   R   T           S      6    ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��    �         -      D                    mosiSignal <= mosiSignal(6 downto 1) & spi_mosi;5�_�   S   U           T      6    ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��    �         -      D                    mosiSignal <= mosiSignal(6 downto 9) & spi_mosi;5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��     �                9                   -- mosiSignal(0)          <= spi_mosi;5�_�   U   Z           V           ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��    �                 5�_�   V   [   Y       Z           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   )   +   +              end process;�   (   *   +                   end if;�   '   )   +                      end if;�   &   (   +      &                  bitCount   <= "000";�   %   '   +                      else �   $   &   +                          end if;�   #   %   +                              �   "   $   +      ,                        bitCount   <= "000";�   !   #   +      =                        ledsData   <= mosiSignal(3 downto 0);�       "   +      1                        outData    <= mosiSignal;�      !   +      4                        spi_miso   <= misoSignal(7);�          +      -                        misoSignal <= inData;�         +      .                    if (bitCount = "111") then�         +      W                    bitCount               <= std_logic_vector(unsigned(bitCount) + 1);�         +      E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);�         +      <                    spi_miso               <= misoSignal(7);�         +      P                    mosiSignal             <= mosiSignal(6 downto 0) & spi_mosi;�         +      "                if (cs = '0') then�         +      $            if rising_edge(clk) then�         +              begin�         +          process (clk)�         +      begin   �         +      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         +      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      '           clk      : in    STD_LOGIC);�   
      +      :           ledsData : out   std_logic_vector (3 downto 0);�   	      +      :           inData   : in    std_logic_vector (7 downto 0);�      
   +      :           outData  : out   std_logic_vector (7 downto 0);�      	   +      &           cs       : in    std_logic;�         +      &           spi_miso : out   STD_LOGIC;�         +      &    Port ( spi_mosi : in    STD_LOGIC;�                D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�                W                    bitCount               <= std_logic_vector(unsigned(bitCount) + 1);�                E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);�                <                    spi_miso               <= misoSignal(7);5�_�   Z   \           [      D    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         +      E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);5�_�   [   ^           \          ����                                                                                                                                                                                                                                                                                                                                         )       v   )    ]��     �         +      K                    misoSignal(7 downto 1) <= misoSignal(6 downto 0) & '0';5�_�   \   _   ]       ^           ����                                                                                                                                                                                                                                                                                                                                                V       ]�     �   )   +   +              end process;�   (   *   +                   end if;�   '   )   +                      end if;�   &   (   +      &                  bitCount   <= "000";�   %   '   +                      else �   $   &   +                          end if;�   #   %   +                              �   "   $   +      ,                        bitCount   <= "000";�   !   #   +      =                        ledsData   <= mosiSignal(3 downto 0);�       "   +      1                        outData    <= mosiSignal;�      !   +      4                        spi_miso   <= misoSignal(7);�          +      -                        misoSignal <= inData;�         +      .                    if (bitCount = "111") then�         +      K                    bitCount   <= std_logic_vector(unsigned(bitCount) + 1);�         +      ?                    misoSignal <= misoSignal(6 downto 0) & '0';�         +      0                    spi_miso   <= misoSignal(7);�         +      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�         +      "                if (cs = '0') then�         +      $            if rising_edge(clk) then�         +              begin�         +          process (clk)�         +      begin   �         +      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         +      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      '           clk      : in    STD_LOGIC);�   
      +      :           ledsData : out   std_logic_vector (3 downto 0);�   	      +      :           inData   : in    std_logic_vector (7 downto 0);�      
   +      :           outData  : out   std_logic_vector (7 downto 0);�      	   +      &           cs       : in    std_logic;�         +      &           spi_miso : out   STD_LOGIC;�         +      &    Port ( spi_mosi : in    STD_LOGIC;�                P                    mosiSignal             <= mosiSignal(6 downto 0) & spi_mosi;�                W                    bitCount               <= std_logic_vector(unsigned(bitCount) + 1);�                ?                    misoSignal <= misoSignal(6 downto 0) & '0';�                <                    spi_miso               <= misoSignal(7);5�_�   ^   `           _          ����                                                                                                                                                                                                                                                                                                                                                V       ]�     �         ,                          �         +    5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                V       ]�    �         ,                          5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                                V       ]�K     �         -             �         ,    5�_�   a   c           b          ����                                                                                                                                                                                                                                                                                                                                                V       ]�g     �         -      K                    bitCount   <= std_logic_vector(unsigned(bitCount) + 1);5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                                V       ]�g     �         -      J                    itCount   <= std_logic_vector(unsigned(bitCount) + 1);5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                V       ]�g     �         -      I                    tCount   <= std_logic_vector(unsigned(bitCount) + 1);5�_�   d   f           e          ����                                                                                                                                                                                                                                                                                                                                                V       ]�h     �         -      H                    Count   <= std_logic_vector(unsigned(bitCount) + 1);5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                                                V       ]�j     �         -      H                    count   <= std_logic_vector(unsigned(bitCount) + 1);5�_�   f   h           g      '    ����                                                                                                                                                                                                                                                                                                                                                V       ]�m     �         -      S                    count   := count +1<= std_logic_vector(unsigned(bitCount) + 1);5�_�   g   i           h           ����                                                                                                                                                                                                                                                                                                                                                  v       ]�p     �      !   -      .                    if (bitCount = "111") then5�_�   h   j           i           ����                                                                                                                                                                                                                                                                                                                                                  v       ]�q     �      !   -      +                    if (Count = "111") then5�_�   i   k           j            ����                                                                                                                                                                                                                                                                                                                                            $       v   $    ]�t     �      !   -      +                    if (count = "111") then5�_�   j   l           k           ����                                                                                                                                                                                                                                                                                                                                            $       v   $    ]�~     �      !   -      '                    if (count = 8) then5�_�   k   m           l           ����                                                                                                                                                                                                                                                                                                                                            $       v   $    ]��     �                 5�_�   l   n           m           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �   *   ,   ,              end process;�   )   +   ,                   end if;�   (   *   ,                      end if;�   '   )   ,      &                  bitCount   <= "000";�   &   (   ,                      else �   %   '   ,                          end if;�   $   &   ,                              �   #   %   ,      ,                        bitCount   <= "000";�   "   $   ,      =                        ledsData   <= mosiSignal(3 downto 0);�   !   #   ,      1                        outData    <= mosiSignal;�       "   ,      4                        spi_miso   <= misoSignal(7);�      !   ,      -                        misoSignal <= inData;�          ,      (                    if (count /= 8) then�         ,      %                    count := count +1�         ,      ?                    misoSignal <= misoSignal(6 downto 0) & '0';�         ,      0                    spi_miso   <= misoSignal(7);�         ,      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�         ,      "                if (cs = '0') then�         ,      $            if rising_edge(clk) then�         ,              begin�         ,      0       variable count: integer range 0 to 8 :=0;�         ,          process (clk)�         ,      begin   �         ,      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         ,      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         ,      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         ,      '           clk      : in    STD_LOGIC);�   
      ,      :           ledsData : out   std_logic_vector (3 downto 0);�   	      ,      :           inData   : in    std_logic_vector (7 downto 0);�      
   ,      :           outData  : out   std_logic_vector (7 downto 0);�      	   ,      &           cs       : in    std_logic;�         ,      &           spi_miso : out   STD_LOGIC;�         ,      &    Port ( spi_mosi : in    STD_LOGIC;�                '                    count   := count +15�_�   m   o           n           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                 5�_�   n   p           o           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;   0                    spi_miso   <= misoSignal(7);   ?                    misoSignal <= misoSignal(6 downto 0) & '0';5�_�   o   r           p          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         (    �         (    5�_�   p   s   q       r          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �          ,                          �          +    5�_�   r   t           s   %       ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �   $   %                                  5�_�   s   u           t           ����                                                                                                                                                                                                                                                                                                                                                  V        ]��     �                D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                  V        ]��     �         *    �         *    5�_�   u   w           v           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                ?                    misoSignal <= misoSignal(6 downto 0) & '0';�                0                    spi_miso   <= misoSignal(7);5�_�   v   x           w           ����                                                                                                                                                                                                                                                                                                                                                V       ]� *     �      !   +    �       !   +    5�_�   w   y           x           ����                                                                                                                                                                                                                                                                                                                                                V       ]� +     �      !          3                       spi_miso   <= misoSignal(7);5�_�   x   z           y   !        ����                                                                                                                                                                                                                                                                                                                            !          %          V       ]� -     �   $   &          ,                        bitCount   <= "000";�   #   %          =                        ledsData   <= mosiSignal(3 downto 0);�   "   $          1                        outData    <= mosiSignal;�   !   #          4                        spi_miso   <= misoSignal(7);�       "          -                        misoSignal <= inData;5�_�   y   {           z   "       ����                                                                                                                                                                                                                                                                                                                            !          %          V       ]� F     �   !   "          0                    spi_miso   <= misoSignal(7);5�_�   z   |           {   $       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ]� W     �   #   %   +      (                    bitCount   <= "000";5�_�   {   }           |   $   "    ����                                                                                                                                                                                                                                                                                                                            $   "       $   &       v   &    ]� Z     �   #   %   +      (                    bitCount   := "000";5�_�   |   ~           }   '        ����                                                                                                                                                                                                                                                                                                                            '   "       '   "       V   "    ]� _     �   &   (   *    �   '   (   *    �   &   '          &                  bitCount   <= "000";5�_�   }              ~   '       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� `     �   &   (          $                    bitCount   := 0;5�_�   ~   �              '       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� a     �   &   (   +      #                   bitCount   := 0;5�_�      �           �   '       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� a     �   &   (   +      "                   itCount   := 0;5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� a     �   &   (   +      !                   tCount   := 0;5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� b     �   &   (   +                          Count   := 0;5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� c     �   #   %   +      $                    bitCount   := 0;5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� c     �   #   %   +      #                    itCount   := 0;5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� c     �   #   %   +      "                    tCount   := 0;5�_�   �   �           �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� d     �   #   %   +      !                    Count   := 0;5�_�   �   �   �       �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� j     �   #   %   +      !                    xount   := 0;5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                            $                     V       ]� m     �   )   +   +              end process;�   (   *   +                   end if;�   '   )   +                      end if;�   &   (   +                          count   := 0;�   %   '   +                      else �   $   &   +                          end if;�   #   %   +      $                    count      := 0;�   "   $   +      9                    ledsData   <= mosiSignal(3 downto 0);�   !   #   +      -                    outData    <= mosiSignal;�       "   +      )                    misoSignal <= inData;�      !   +      0                    spi_miso   <= misoSignal(7);�          +                       else�         +      B                       misoSignal <= misoSignal(6 downto 0) & '0';�         +      3                       spi_miso   <= misoSignal(7);�         +      (                    if (count /= 8) then�         +      %                    count := count +1�         +      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�         +      "                if (cs = '0') then�         +      $            if rising_edge(clk) then�         +              begin�         +      0       variable count: integer range 0 to 8 :=0;�         +          process (clk)�         +      begin   �         +      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         +      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      '           clk      : in    STD_LOGIC);�   
      +      :           ledsData : out   std_logic_vector (3 downto 0);�   	      +      :           inData   : in    std_logic_vector (7 downto 0);�      
   +      :           outData  : out   std_logic_vector (7 downto 0);�      	   +      &           cs       : in    std_logic;�         +      &           spi_miso : out   STD_LOGIC;�         +      &    Port ( spi_mosi : in    STD_LOGIC;�      !          0                    spi_miso   <= misoSignal(7);�   #   %          !                    count   := 0;�   "   $          9                    ledsData   <= mosiSignal(3 downto 0);�   !   #          -                    outData    <= mosiSignal;�       "          )                    misoSignal <= inData;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]� z    �   )   +   +              end process;�   (   *   +                   end if;�   '   )   +                      end if;�   &   (   +                          count   := 0;�   %   '   +                      else �   $   &   +                          end if;�   #   %   +      $                    count      := 0;�   "   $   +      9                    ledsData   <= mosiSignal(3 downto 0);�   !   #   +      -                    outData    <= mosiSignal;�       "   +      )                    misoSignal <= inData;�      !   +      0                    spi_miso   <= misoSignal(7);�          +                       else�         +      B                       misoSignal <= misoSignal(6 downto 0) & '0';�         +      3                       spi_miso   <= misoSignal(7);�         +      (                    if (count /= 8) then�         +      *                    count      := count +1�         +      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�         +      "                if (cs = '0') then�         +      $            if rising_edge(clk) then�         +              begin�         +      0       variable count: integer range 0 to 8 :=0;�         +          process (clk)�         +      begin   �         +      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         +      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      '           clk      : in    STD_LOGIC);�   
      +      :           ledsData : out   std_logic_vector (3 downto 0);�   	      +      :           inData   : in    std_logic_vector (7 downto 0);�      
   +      :           outData  : out   std_logic_vector (7 downto 0);�      	   +      &           cs       : in    std_logic;�         +      &           spi_miso : out   STD_LOGIC;�         +      &    Port ( spi_mosi : in    STD_LOGIC;�                D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�                %                    count := count +15�_�   �   �           �      *    ����                                                                                                                                                                                                                                                                                                                                                V       ]� �    �         +      *                    count      := count +15�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                               !       %          V   !    ]�&    �   #   %          $                    count      := 0;�   "   $          9                    ledsData   <= mosiSignal(3 downto 0);�   !   #          -                    outData    <= mosiSignal;�       "          )                    misoSignal <= inData;�      !          0                    spi_miso   <= misoSignal(7);�                                  else5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]�&%    �   )   +   +              end process;�   (   *   +                   end if;�   '   )   +                      end if;�   &   (   +                         count := 0;�   %   '   +                      else �   $   &   +                          end if;�   #   %   +      '                       count      := 0;�   "   $   +      <                       ledsData   <= mosiSignal(3 downto 0);�   !   #   +      0                       outData    <= mosiSignal;�       "   +      ,                       misoSignal <= inData;�      !   +      3                       spi_miso   <= misoSignal(7);�          +                          else�         +      B                       misoSignal <= misoSignal(6 downto 0) & '0';�         +      3                       spi_miso   <= misoSignal(7);�         +      (                    if (count /= 8) then�         +      +                    count      := count +1;�         +      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�         +      "                if (cs = '0') then�         +      $            if rising_edge(clk) then�         +              begin�         +      0       variable count: integer range 0 to 8 :=0;�         +          process (clk)�         +      begin   �         +      I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');�         +      I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');�         +      '           clk      : in    STD_LOGIC);�   
      +      :           ledsData : out   std_logic_vector (3 downto 0);�   	      +      :           inData   : in    std_logic_vector (7 downto 0);�      
   +      :           outData  : out   std_logic_vector (7 downto 0);�      	   +      &           cs       : in    std_logic;�         +      &           spi_miso : out   STD_LOGIC;�         +      &    Port ( spi_mosi : in    STD_LOGIC;�   &   (                              count   := 0;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�&�     �                3                       spi_miso   <= misoSignal(7);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�&�     �         *    �         *    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                V       ]�&�     �                3                       spi_miso   <= misoSignal(7);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�&�    �                 3                       spi_miso   <= misoSignal(7);5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/p     �                I    signal bitCount   : std_logic_vector (2 downto 0) := (others => '0');5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/�     �         )      (                    if (count /= 8) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/�    �         )      (                    if (count <= 8) then5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/�    �         )      '                    if (count < 8) then5�_�   �   �           �      *    ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/�     �         )      0       variable count: integer range 0 to 8 :=0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�/�   ! �         )      (                    if (count <= 8) then5�_�   �   �           �       %    ����                                                                                                                                                                                                                                                                                                                                %           .       v   .    ]�0v     �      !   )      0                       outData    <= mosiSignal;�       !   )    5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   .       v   .    ]�0�     �       "   )      <                       ledsData   <= mosiSignal(3 downto 0);�   !   "   )    5�_�   �   �           �   !   F    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�     �       "   )      S                       ledsData   <= mosiSignal(6 downto 0) & spi_mosi(3 downto 0);5�_�   �   �           �   !   G    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�     �       "   )      U                       ledsData   <= mosiSignal(6 downto 0) & spi_mosi)h(3 downto 0);5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�   " �       "   )      T                       ledsData   <= mosiSignal(6 downto 0) & spi_mosi)(3 downto 0);5�_�   �   �           �   !   G    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�     �       "   )      U                       ledsData   <= (mosiSignal(6 downto 0) & spi_mosi)(3 downto 0);5�_�   �   �           �   !   1    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�     �       "   )      T                       ledsData   <= (mosiSignal(6 downto 0) & spi_mosi(3 downto 0);5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   E       v   .    ]�0�     �       "   )      T                       ledsData   <= (mosiSignal(2 downto 0) & spi_mosi(3 downto 0);5�_�   �   �           �   !   F    ����                                                                                                                                                                                                                                                                                                                            !   F       !   Q       v   Q    ]�0�   # �       "   )      S                       ledsData   <= mosiSignal(2 downto 0) & spi_mosi(3 downto 0);5�_�   �   �           �      *    ����                                                                                                                                                                                                                                                                                                                            !   F       !   Q       v   Q    ]�0�   ( �         )      0       variable count: integer range 0 to 9 :=0;5�_�   �   �   �       �   
        ����                                                                                                                                                                                                                                                                                                                               /          /       V   /    ]�2�   ) �   	             :           inData   : in    std_logic_vector (7 downto 0);5�_�   �   �           �   
   9    ����                                                                                                                                                                                                                                                                                                                                                             ]���   + �   	      )      :           inData   : in    std_logic_vector (7 downto 0),5�_�   �               �      %    ����                                                                                                                                                                                                                                                                                                                                                             ]���     �         )      -                 spi_miso   <= misoSignal(7);   (                 count      := count +1;5�_�   �   �   �   �   �           ����                                                                                                                                                                                                                                                                                                                               /          /       V   /    ]�2W     �              5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                               /          /       V   /    ]�2X     �         (    �         (      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   �   �       �   �       /    ����                                                                                                                                                                                                                                                                                                                            !   F       !   Q       v   Q    ]�2;     �      !   )      J                       outData    <= mosiSignal;--(6 downto 0) & spi_mosi;5�_�   �               �       0    ����                                                                                                                                                                                                                                                                                                                            !   F       !   Q       v   Q    ]�2?   % �      !   )      K                       outData    <= mosiSignal; --(6 downto 0) & spi_mosi;5�_�   �   �       �   �           ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�'�     �              5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�'�     �         )    �         )      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                               "          "       V   "    ]�'�     �                G                       mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                            !   %       !   =       v   =    ]�'�     �   !   "   *    �       !   *      G                       mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   =       v   =    ]�'�    �       "   +      .                       mosiSignal <= spi_mosi;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   =       v   =    ]�'�     �       "   +      ?                       mosiSignal <= others => '0') & spi_mosi;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   3       v   3    ]�'�    �       "   +      @                       mosiSignal <= (others => '0') & spi_mosi;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   %       !   3       v   3    ]�(     �       "   +      ?                       mosiSignal <= others => '0') & spi_mosi;5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                            !   .       !   ;       v   ;    ]�(     �       "   +      H                       mosiSignal <= "0000000"others => '0') & spi_mosi;5�_�   �               �   !   .    ����                                                                                                                                                                                                                                                                                                                            !   .       !   ;       v   ;    ]�(    �       "   +      :                       mosiSignal <= "0000000" & spi_mosi;5�_�   �           �   �   $       ����                                                                                                                                                                                                                                                                                                                            '           '   #       V   "    ]� f     �   #   %   +                             := 0;5�_�   p           r   q          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         +    �         +      D                    mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;   0                    spi_miso   <= misoSignal(7);   ?                    misoSignal <= misoSignal(6 downto 0) & '0';5�_�   \           ^   ]           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         +      Peeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   <eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ?eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Weeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   V       X   Z   Y           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         +      Deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   <eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Weeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   V       W   Y   X           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         +      Deeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   <eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Weeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   V           X   W           ����                                                                                                                                                                                                                                                                                                                                         <       V   <    ]��     �                C                   mosiSignal <= mosiSignal(6 downto 0) & spi_mosi;�                ;                   spi_miso               <= misoSignal(7);�                D                   misoSignal(7 downto 1) <= misoSignal(6 downto 0);�                V                   bitCount               <= std_logic_vector(unsigned(bitCount) + 1);5�_�   >           @   ?          ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         ,      Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   .eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   .eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   Ieeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5��