Vim�UnDo� �>��˷)R���x�<�{���G:l�C��   ?                 Z  Z  Z  Z  Y    ^Y   � _�                            ����                                                                                                                                                                                                                                                                                                                                                             ]��     �               entity negador_tb is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]��     �               !architecture arq of negador_tb is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             ]��"     �      	            component negador is5�_�                    	        ����                                                                                                                                                                                                                                                                                                                            	          	          V       ]��%     �      
               generic(            N: std_logic := '1'5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	          	          V       ]��&     �      	          "      generic( N: std_logic := '1'5�_�                    	       ����                                                                                                                                                                                                                                                                                                                            	          	          V       ]��'     �      	                );5�_�                            ����                                                                                                                                                                                                                                                                                                                            	          	          V       ]��-     �      X       5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                       *           V        ]��2     �             $   R----------------------------------------------------------------------------------   -- Company:    -- Engineer:    --    &-- Create Date: 12/04/2019 04:59:29 PM   -- Design Name:    #-- Module Name: spi28b - Behavioral   -- Project Name:    -- Target Devices:    -- Tool Versions:    -- Description:    --    -- Dependencies:    --    -- Revision:   -- Revision 0.01 - File Created   -- Additional Comments:   --    R----------------------------------------------------------------------------------           library IEEE;   use IEEE.STD_LOGIC_1164.ALL;   use IEEE.numeric_std.all;    use IEEE.std_logic_unsigned.all;       7-- Uncomment the following library declaration if using   6-- arithmetic functions with Signed or Unsigned values   --use IEEE.NUMERIC_STD.ALL;       ?-- Uncomment the following library declaration if instantiating   &-- any Xilinx leaf cells in this code.   --library UNISIM;   --use UNISIM.VComponents.all;       entity spi28b is5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                                                V       ]��6     �                &    Port ( spi_mosi : in    STD_LOGIC;   &           spi_miso : out   STD_LOGIC;   &           cs       : in    std_logic;   :           outData  : out   std_logic_vector (7 downto 0);   :           inData   : in    std_logic_vector (7 downto 0);   :           ledsData : out   std_logic_vector (3 downto 0);   '           clk      : in    STD_LOGIC);   end spi28b;5�_�   	              
   .        ����                                                                                                                                                                                                                                                                                                                                                V       ]��:     �   -   6   A    �   .   /   A    5�_�   
                 4   %    ����                                                                                                                                                                                                                                                                                                                                                V       ]��>     �   3   6   I      '           clk      : in    STD_LOGIC);5�_�                    6        ����                                                                                                                                                                                                                                                                                                                                                V       ]��A     �   5   6          end spi28b;5�_�                    6        ����                                                                                                                                                                                                                                                                                                                            6          ;          V       ]��C     �   5   6                port(            a:   in  std_logic;            b:   out std_logic;            rst: in  std_logic;            clk: in  std_logic         );5�_�                    6       ����                                                                                                                                                                                                                                                                                                                            6          6          V       ]��D     �   6   8   C    5�_�                    8        ����                                                                                                                                                                                                                                                                                                                            8          ;          V       ]��G     �   7   8          $   signal a_tb:    std_logic := '0';      signal b_tb:    std_logic;   $   signal clk_tb:  std_logic := '0';      signal rst_tb:  std_logic;5�_�                    9        ����                                                                                                                                                                                                                                                                                                                            9           <           V        ]��I     �   8   9          %   a_tb   <= not a_tb   after 200 ns;   $   clk_tb <= not clk_tb after 20 ns;      rst_tb <= '0';    5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            9           9           V        ]��M     �   8   :   <         aa: negador5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            9           9           V        ]��P     �   8   :   <         spi_inst: negador5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            9           9           V        ]��V     �   9   :                generic map(N=>'0')5�_�                    .       ����                                                                                                                                                                                                                                                                                                                            9           9           V        ]��Z     �   -   /   ;      &    Port ( spi_mosi : in    STD_LOGIC;5�_�                   :        ����                                                                                                                                                                                                                                                                                                                            :           :           V        ]��e     �   9   ;   ;    �   :   ;   ;    5�_�                    :        ����                                                                                                                                                                                                                                                                                                                            :          :          V       ]��j     �   9   B   ;    �   :   ;   ;    �   9   :          ;      port map(a=>a_tb, b=>b_tb, clk=>clk_tb, rst=>rst_tb);5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            :           A   	       V       ]��o     �   9   ;   C      &    port ( spi_mosi : in    STD_LOGIC;5�_�                   :        ����                                                                                                                                                                                                                                                                                                                            :   )       A   	       V   	    ]�Ƀ     �   @   B          
        );�   >   @          :           ledsData : out   std_logic_vector (3 downto 0);�   =   ?          :           inData   : in    std_logic_vector (7 downto 0);�   <   >          :           outData  : out   std_logic_vector (7 downto 0);�   ;   =          &           cs       : in    std_logic;�   :   <          &           spi_miso : out   STD_LOGIC;�   9   ;          *    port map ( spi_mosi : in    STD_LOGIC;5�_�                    A   	    ����                                                                                                                                                                                                                                                                                                                            :   )       A   	       V   	    ]�Ɇ     �   @   B   C      
        ),5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            ;          @                 ]�ɗ     �   ;   A   C      &           cs       : in    std_logic,   :           outData  : out   std_logic_vector (7 downto 0),   :           inData   : in    std_logic_vector (7 downto 0),   :           ledsData : out   std_logic_vector (3 downto 0),   %           clk      : in    STD_LOGIC�   :   <   C      &           spi_miso : out   STD_LOGIC,5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            ;          @                 ]�ɥ     �   :   B   C      (           spi_miso =>  out   STD_LOGIC,   (           cs       =>  in    std_logic,   <           outData  =>  out   std_logic_vector (7 downto 0),   <           inData   =>  in    std_logic_vector (7 downto 0),   <           ledsData =>  out   std_logic_vector (3 downto 0),   '           clk      =>  in    STD_LOGIC   
        );�   ;   <   C    �   :   A   C      )           spi_miso => : out   STD_LOGIC,   )           cs       => : in    std_logic,   =           outData  => : out   std_logic_vector (7 downto 0),   =           inData   => : in    std_logic_vector (7 downto 0),   =           ledsData => : out   std_logic_vector (3 downto 0),   (           clk      => : in    STD_LOGIC5�_�                    ;        ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]�ɫ     �   :   <   C                  spi_miso => spi_miso �   :   A   C      1           spi_miso => spi_miso  out   STD_LOGIC,   1           cs       => cs        in    std_logic,   E           outData  => outData   out   std_logic_vector (7 downto 0),   E           inData   => inData    in    std_logic_vector (7 downto 0),   E           ledsData => ledsData  out   std_logic_vector (3 downto 0),   0           clk      => clk       in    STD_LOGIC5�_�                     @        ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]�ɲ     �   ?   A   C      !           clk      => clk      ,5�_�      !               @       ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]�ɳ     �   ?   A   C                  clk      => clk      5�_�       "           !   B       ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]�ɶ     �   A   B          ;      port map(a=>a_tb, b=>b_tb, clk=>clk_tb, rst=>rst_tb);5�_�   !   #           "   :       ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]�ɽ     �   9   ;   B      *    port map ( spi_mosi : in    STD_LOGIC,5�_�   "   $           #   :       ����                                                                                                                                                                                                                                                                                                                            ;           @   0       ���    ]���     �   9   ;   B      -    port map ( spi_mosi => : in    STD_LOGIC,5�_�   #   %           $   :       ����                                                                                                                                                                                                                                                                                                                            :          :          v       ]���     �   9   ;   B      ,    port map ( spi_mosi =>  in    STD_LOGIC,�   :   ;   B    5�_�   $   &           %   :   #    ����                                                                                                                                                                                                                                                                                                                            :          :          v       ]���     �   9   ;   B      4    port map ( spi_mosi => spi_mosi in    STD_LOGIC,5�_�   %   '           &   ;       ����                                                                                                                                                                                                                                                                                                                            ;          @                 ]���     �   ;   A   B      !           cs       => cs       ,   !           outData  => outData  ,   !           inData   => inData   ,   !           ledsData => ledsData ,              clk      => clk�   :   <   B      !           spi_miso => spi_miso ,5�_�   &   )           '   :   #    ����                                                                                                                                                                                                                                                                                                                            ;          @                 ]���     �   9   ;   B      $    port map ( spi_mosi => spi_mosi,5�_�   '   *   (       )   :   #    ����                                                                                                                                                                                                                                                                                                                            :   #       ?   #          #    ]���     �   9   ;   B      %    port map ( spi_mosi => spi_mosi ,5�_�   )   +           *   ;   #    ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   :   <   B      %           spi_miso     => spi_miso ,�   ;   <   B    5�_�   *   ,           +   <       ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   ;   =   B      %           cs           => cs       ,�   <   =   B    5�_�   +   -           ,   =   "    ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   <   >   B      %           outData      => outData  ,�   =   >   B    5�_�   ,   .           -   >   !    ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   =   ?   B      %           inData       => inData   ,�   >   ?   B    5�_�   -   /           .   ?   #    ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   >   @   B      %           ledsData     => ledsData ,�   ?   @   B    5�_�   .   0           /   @       ����                                                                                                                                                                                                                                                                                                                            :   #       :   %       v   %    ]���     �   ?   A   B                 clk          => clk�   @   A   B    5�_�   /   1           0           ����                                                                                                                                                                                                                                                                                                                                       )          V        ]��     �             "   $architecture Behavioral of spi28b is   I    signal mosiSignal : std_logic_vector (7 downto 0) := (others => '0');   I    signal misoSignal : std_logic_vector (7 downto 0) := (others => '0');   D    signal bitCount   : std_logic_vector (7 downto 0) := "00000001";       begin          process (clk)               begin   $            if rising_edge(clk) then   "                if (cs = '0') then                                                E                    mosiSignal(7 downto 1) <= mosiSignal(6 downto 0);   .                    mosiSignal(0) <= spi_mosi;                          .                    spi_miso <= misoSignal(7);   E                    misoSignal(7 downto 1) <= misoSignal(6 downto 0);                          A                    bitCount(7 downto 1) <= bitCount(6 downto 0);       3                    if (bitCount = "00000000") then   -                        misoSignal <= inData;   4                        spi_miso   <= misoSignal(7);   1                        outData    <= mosiSignal;   =                        ledsData   <= mosiSignal(3 downto 0);   0                        bitCount   <="00000001";                                                  end if;                   else    *                  bitCount   <="00000001";                   end if;                end if;           end process;5�_�   0   2           1           ����                                                                                                                                                                                                                                                                                                                                                  V        ]��
     �                     5�_�   1   3           2           ����                                                                                                                                                                                                                                                                                                                                                  V        ]��    �                end Behavioral;5�_�   2   4           3           ����                                                                                                                                                                                                                                                                                                                                                             ]���     �                5�_�   3   5           4           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �             �             5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                       ]��     �         %          spi_mosi_tb ,�         %      (    port map ( spi_mosi => spi_mosi_tb ,   (           spi_miso     => spi_miso_tb ,   (           cs           => cs_tb       ,   (           outData      => outData_tb  ,   (           inData       => inData_tb   ,   (           ledsData     => ledsData_tb ,   !           clk          => clk_tb5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                       ]��     �         %          signal spi_mosi_tb        signal spi_miso_tb        signal cs_tb              signal outData_tb         signal inData_tb          signal ledsData_tb        signal clk_tb    �         %    �         %          signal spi_mosi_tb ,       signal spi_miso_tb ,       signal cs_tb       ,       signal outData_tb  ,       signal inData_tb   ,       signal ledsData_tb ,5�_�   6   :           7      (    ����                                                                                                                                                                                                                                                                                                                                         <              ]��(    �         %      (    signal clk_tb      : in    STD_LOGIC5�_�   7   ;   8       :          ����                                                                                                                                                                                                                                                                                                                                                       ]�ˌ    �         %      )    signal spi_mosi_tb : in    STD_LOGIC;   )    signal spi_miso_tb : out   STD_LOGIC;   )    signal cs_tb       : in    std_logic;   =    signal outData_tb  : out   std_logic_vector (7 downto 0);   =    signal inData_tb   : in    std_logic_vector (7 downto 0);   =    signal ledsData_tb : out   std_logic_vector (3 downto 0);   )    signal clk_tb      : in    STD_LOGIC;5�_�   :   <           ;           ����                                                                                                                                                                                                                                                                                                                                                             ]���     �         %    �         %    5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             ]���     �          (    5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                             ]���     �         )    �         )    5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                             ]���     �         *      #    signal clk_tb      : STD_LOGIC;5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             ]���    �                %   a_tb   <= not a_tb   after 200 ns;5�_�   ?   A           @   !   &    ����                                                                                                                                                                                                                                                                                                                            !   &       &   &          &    ]��7    �       '   )      (    port map ( spi_mosi => spi_mosi_tb ,   (           spi_miso     => spi_miso_tb ,   (           cs           => cs_tb       ,   (           outData      => outData_tb  ,   (           inData       => inData_tb   ,   (           ledsData     => ledsData_tb ,5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                            !   &       &   &          &    ]��d     �         )    5�_�   A   C           B   )       ����                                                                                                                                                                                                                                                                                                                            "   &       '   &          &    ]��i   
 �   )   +   *    5�_�   B   D           C   !       ����                                                                                                                                                                                                                                                                                                                                                             ]��     �       "   +         spi_inst: spi5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                             ]��    �      	   +         component spi is5�_�   D   F           E      "    ����                                                                                                                                                                                                                                                                                                                                                             ]��b    �         +      #    signal clk_tb      : STD_LOGIC;5�_�   E   G           F            ����                                                                                                                                                                                                                                                                                                                                                             ]���    �       #   ,         �       "   +    5�_�   F   H           G   !        ����                                                                                                                                                                                                                                                                                                                                                             ]���     �       -   -       5�_�   G   I           H   !        ����                                                                                                                                                                                                                                                                                                                                                             ]��     �       "   8      VECTOR <= "00000000";5�_�   H   J           I   !       ����                                                                                                                                                                                                                                                                                                                                                             ]��     �       "   8         VECTOR <= "00000000";5�_�   I   K           J   !       ����                                                                                                                                                                                                                                                                                                                                                             ]��     �       "   8         data_out <= "00000000";5�_�   J   L           K   !       ����                                                                                                                                                                                                                                                                                                                                                             ]��     �       "   8         data_in <= "00000000";5�_�   K   M           L   !       ����                                                                                                                                                                                                                                                                                                                                                             ]��'     �       "   8         data_in <= "00000001";5�_�   L   N           M   #       ����                                                                                                                                                                                                                                                                                                                                                             ]��0     �   "   $   8      	for i in 0 to 255 loop5�_�   M   O           N   $       ����                                                                                                                                                                                                                                                                                                                            $          $   	       v       ]��6     �   #   %   8      		WAIT FOR period;5�_�   N   P           O   $       ����                                                                                                                                                                                                                                                                                                                            $          $   	       v       ]��8     �   #   %   8      		WAIT FOR period;5�_�   O   Q           P   $       ����                                                                                                                                                                                                                                                                                                                            $          $   	       v       ]��<     �   #   %   8      		wait for period;5�_�   P   R           Q   %       ����                                                                                                                                                                                                                                                                                                                            %          %          v       ]��P     �   $   &   8      6		VECTOR <= STD_LOGIC_VECTOR (unsigned(VECTOR) + '1');5�_�   Q   S           R   %       ����                                                                                                                                                                                                                                                                                                                            %          %          v       ]��R     �   $   &   8      6		vector <= STD_LOGIC_VECTOR (unsigned(VECTOR) + '1');5�_�   R   T           S   %   *    ����                                                                                                                                                                                                                                                                                                                            %          %          v       ]��Y     �   $   &   8      9		inData_tb <= STD_LOGIC_VECTOR (unsigned(VECTOR) + '1');5�_�   S   U           T   %       ����                                                                                                                                                                                                                                                                                                                            %          %          v   "    ]��a     �   $   &   8      <		inData_tb <= STD_LOGIC_VECTOR (unsigned(inData_tb) + '1');5�_�   T   V           U   &       ����                                                                                                                                                                                                                                                                                                                            %          %          v   "    ]��c     �   %   &          		5�_�   U   W           V   &       ����                                                                                                                                                                                                                                                                                                                            %          %          v   "    ]��h     �   %   &          		WAIT FOR period;5�_�   V   X           W   &       ����                                                                                                                                                                                                                                                                                                                            &          &          v   
    ]��l     �   %   '   6      
	END LOOP;5�_�   W   Y           X   (       ����                                                                                                                                                                                                                                                                                                                            &          &          v   
    ]��z     �   '   (          	wait FOR period;5�_�   X   Z           Y   (        ����                                                                                                                                                                                                                                                                                                                            &          &          v   
    ]��z     �   '   (           5�_�   Y   [           Z   (        ����                                                                                                                                                                                                                                                                                                                            &          &          v   
    ]��{     �   '   (           5�_�   Z   \           [            ����                                                                                                                                                                                                                                                                                                                            &          &          v   
    ]��     �                  5�_�   [   ]           \   !        ����                                                                                                                                                                                                                                                                                                                            %          %          v   
    ]��     �       $   2       5�_�   \   ^           ]   $        ����                                                                                                                                                                                                                                                                                                                            $          '          V       ]��     �   #   (   4      	for i in 0 to 10 loop   		wait for 100ns;   <		inData_tb <= std_logic_vector (unsigned(inData_tb) + '1');   
	end loop;5�_�   ]   _           ^   '       ����                                                                                                                                                                                                                                                                                                                            $          '          V       ]��     �   '   )   4    �   '   (   4    5�_�   ^   `           _   '       ����                                                                                                                                                                                                                                                                                                                            $          '          V       ]���     �   '   )   6            �   '   )   5    5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                 V       ]���    �   3   5   6      
        );�   2   4   6      !           clk          => clk_tb�   1   3   6      '           ledsData     => ledsData_tb,�   0   2   6      '           inData       => inData_tb  ,�   /   1   6      '           outData      => outData_tb ,�   .   0   6      '           cs           => cs_tb      ,�   -   /   6      '           spi_miso     => spi_miso_tb,�   ,   .   6      '    port map ( spi_mosi => spi_mosi_tb,�   +   -   6         spi_inst: spi28b�   )   +   6      	�   '   )   6         end process;�   &   (   6            end loop;�   %   '   6      C         inData_tb <= std_logic_vector (unsigned(inData_tb) + '1');�   $   &   6               wait for 100ns;�   #   %   6            for i in 0 to 10 loop�   "   $   6         begin�   !   #   6         loop_proc: process�      !   6         inData_tb <= "00000001";�          6         rst_tb    <= '0';�         6      '   clk_tb    <= not clk_tb after 20 ns;�         6            �         6      #    signal rst_tb      : STD_LOGIC;�         6      *    signal clk_tb      : STD_LOGIC := '0';�         6      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         6      7    signal inData_tb   : std_logic_vector (7 downto 0);�         6      7    signal outData_tb  : std_logic_vector (7 downto 0);�         6      #    signal cs_tb       : std_logic;�         6      #    signal spi_miso_tb : STD_LOGIC;�         6      #    signal spi_mosi_tb : STD_LOGIC;�         6         end component;�         6      
        );�         6      %           clk      : in    STD_LOGIC�         6      :           ledsData : out   std_logic_vector (3 downto 0);�         6      :           inData   : in    std_logic_vector (7 downto 0);�         6      :           outData  : out   std_logic_vector (7 downto 0);�   
      6      &           cs       : in    std_logic;�   	      6      &           spi_miso : out   STD_LOGIC;�      
   6      &    port ( spi_mosi : in    STD_LOGIC;�      	   6         component spi28b is�                $   clk_tb <= not clk_tb after 20 ns;�      !             inData_tb <= "00000001";�                    rst_tb <= '0';5�_�   `   b           a   )        ����                                                                                                                                                                                                                                                                                                                            )           *           V        ]���    �   (   )                 5�_�   a   c           b           ����                                                                                                                                                                                                                                                                                                                            )           )           V        ]���    �                 5�_�   b   d           c   $       ����                                                                                                                                                                                                                                                                                                                            (           (           V        ]���    �   #   %   3               wait for 100ns;5�_�   c   e           d           ����                                                                                                                                                                                                                                                                                                                            (           (           V        ]��     �         3    �         3    5�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                            )           )           V        ]��     �                 5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                            (           (           V        ]��    �         3    5�_�   f   h           g   "       ����                                                                                                                                                                                                                                                                                                                            )           )           V        ]��'     �   "   $   5            �   "   $   4    5�_�   g   i           h   #        ����                                                                                                                                                                                                                                                                                                                            #          #          V       ]��@     �   "   #                variable i: integer := 0;5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                            #          #          V       ]��B     �         4    �         4    5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]��C     �         5            variable i: integer := 0;5�_�   j   l           k          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]��D    �         5           variable i: integer := 0;5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                            $          $          V       ]��^     �         5    �         5    5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                            %          %          V       ]��`    �         6      use ieee.std_logic_1164.all;5�_�   m   o           n           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                    variable i: integer := 0;5�_�   n   p           o   $       ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �   #   %   5    �   $   %   5    5�_�   o   q           p           ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �                use ieee.std_logic_arith.all;5�_�   p   r           q   '   >    ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �   &   (   5      C         inData_tb <= std_logic_vector (unsigned(inData_tb) + '1');5�_�   q   s           r   '   ?    ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �   &   (   5      B         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1');5�_�   r   t           s      6    ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �         5      7    signal inData_tb   : std_logic_vector (7 downto 0);5�_�   s   u           t      :    ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �         5      E    signal inData_tb   : std_logic_vector (7 downto 0) := '00000000';5�_�   t   v           u      C    ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �         5      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000';5�_�   u   w           v           ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �                    inData_tb <= "00000001";5�_�   v   x           w   "        ����                                                                                                                                                                                                                                                                                                                                                V       ]��I     �   !   #   4          variable i: integer := 0;5�_�   w   y           x           ����                                                                                                                                                                                                                                                                                                                                                V       ]��J     �          4    �          4    5�_�   x   z           y           ����                                                                                                                                                                                                                                                                                                                                                V       ]��M     �      !   5         rst_tb    <= '0';5�_�   y   {           z           ����                                                                                                                                                                                                                                                                                                                                                V       ]��R    �      !   5         cs_tb    <= '0';5�_�   z   |           {      "    ����                                                                                                                                                                                                                                                                                                                                                V       ]��     �         5      #    signal cs_tb       : std_logic;5�_�   {   }           |           ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �      !   5         cs_tb    <= '0' after 60 ns;5�_�   |   ~           }           ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �      !   5         cs_tb    <= '1' after 60 ns;5�_�   }              ~      '    ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �         5      *    signal clk_tb      : STD_LOGIC := '0';5�_�   ~   �                 '    ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �         5      *    signal clk_tb      : STD_LOGIC := '1';5�_�      �           �      '    ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �         5      *    signal cs_tb       : std_logic := '0';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                V       ]���     �         5      *    signal cs_tb       : std_logic := '2';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                V       ]���    �         5      *    signal clk_tb      : STD_LOGIC := '1';5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]��    �   %   '   5               wait for 100 ns;5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                V       ]��,     �          5         rst_tb    <= '0';5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                V       ]��,     �         5      '   clk_tb    <= not clk_tb after 20 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�=     �   %   '   5               wait for 1000 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�>     �   %   '   5               wait for 8000 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�>     �   %   '   5               wait for 800 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�D     �   %   '   5               wait for 80 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�E     �   %   '   5               wait for 16080 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]�F     �   %   '   5               wait for 1600 ns;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�L   ! �      !   5         cs_tb    <= '0' after 60 ns;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ]�e   " �      !   5         cs_tb    <= '0' after 0 ns;5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                V       ]��   # �   %   '   5               wait for 160 ns;5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                                                V       ]�5     �   )   ,   6         �   )   +   5    5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�<     �   *   3   7    �   +   ,   7    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�?     �   *   ,   ?         loop_proc: process5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�D     �   *   ,   ?         spioop_proc: process5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�D     �   *   ,   ?         spiop_proc: process5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�D     �   *   ,   ?         spip_proc: process5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�F     �   *   ,   ?         spi_proc: process5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�I     �   +   .   @            �   +   -   ?    5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]�r     �   ,   /   A               spi_mosi_tb <=5�_�   �   �           �   -   $    ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]��     �   ,   .   B      $         spi_mosi_tb <= inData_tb(7)5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]��     �   .   0   B    5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]��     �   -   /   C       5�_�   �   �   �       �   .        ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]��     �   .   0   D      	         �   .   0   C    5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��     �   0   2   D         variable i: integer := 0;      begin5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            1          5          V       ]��     �   0   1          "   variable i: integer := 0; begin         for i in 0 to 10 loop            wait for 320 ns;   A         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);         end loop;5�_�   �   �           �   0        ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��   $ �   /   0           5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            0          0          V       ]��   % �   +   -   >            �   +   -   =    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��     �   *   ,   >         spi_proc: process(clk)5�_�   �   �   �       �   -       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��   & �   ,   .   >            if(rising_edge(clk)) then5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            /   !       .   !       V   !    ]�   ' �   ;   =   >      
        );�   :   <   >      !           clk          => clk_tb�   9   ;   >      '           ledsData     => ledsData_tb,�   8   :   >      '           inData       => inData_tb  ,�   7   9   >      '           outData      => outData_tb ,�   6   8   >      '           cs           => cs_tb      ,�   5   7   >      '           spi_miso     => spi_miso_tb,�   4   6   >      '    port map ( spi_mosi => spi_mosi_tb,�   3   5   >         spi_inst: spi28b�   0   2   >         end process;�   /   1   >            end if;�   .   0   >      4         inData_tb   <= inData_tb(6 downto 1) & '0';�   -   /   >      %         spi_mosi_tb <= inData_tb(7);�   ,   .   >      "      if(rising_edge(clk_tb)) then�   +   -   >         begin�   *   ,   >         spi_proc: process(clk_tb)�   (   *   >         end process;�   '   )   >            end loop;�   &   (   >      A         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);�   %   '   >               wait for 320 ns;�   $   &   >            for i in 0 to 10 loop�   #   %   >         begin�   "   $   >         variable i: integer := 0;�   !   #   >         loop_proc: process�      !   >         cs_tb    <= '0' after 1 ns;�          >         rst_tb   <= '0';�         >      &   clk_tb   <= not clk_tb after 20 ns;�         >            �         >      #    signal rst_tb      : STD_LOGIC;�         >      *    signal clk_tb      : STD_LOGIC := '0';�         >      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         >      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         >      7    signal outData_tb  : std_logic_vector (7 downto 0);�         >      *    signal cs_tb       : std_logic := '1';�         >      #    signal spi_miso_tb : STD_LOGIC;�         >      #    signal spi_mosi_tb : STD_LOGIC;�         >         end component;�         >      
        );�         >      %           clk      : in    STD_LOGIC�         >      :           ledsData : out   std_logic_vector (3 downto 0);�         >      :           inData   : in    std_logic_vector (7 downto 0);�         >      :           outData  : out   std_logic_vector (7 downto 0);�         >      &           cs       : in    std_logic;�   
      >      &           spi_miso : out   STD_LOGIC;�   	      >      &    port ( spi_mosi : in    STD_LOGIC;�      
   >         component spi28b is�   -   /          %         spi_mosi_tb <= inData_tb(7);�   .   0          2         inData_tb <= inData_tb(6 downto 1) & '0';5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            /   !       .   !       V   !    ]�      �   ,   .   >      "      if(rising_edge(clk_tb)) then5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                            /   !       .   !       V   !    ]�!   ( �   ,   .   >      "      if rising_edge(clk_tb)) then5�_�   �   �           �   /   +    ����                                                                                                                                                                                                                                                                                                                            /   !       .   !       V   !    ]�'   ) �   .   0   >      4         inData_tb   <= inData_tb(6 downto 1) & '0';5�_�   �   �           �   +   	    ����                                                                                                                                                                                                                                                                                                                            /   !       .   !       V   !    ]��     �   +   -   >    �   +   ,   >    5�_�   �   �           �   ,        ����                                                                                                                                                                                                                                                                                                                            0   !       /   !       V   !    ]��     �   +   .   ?       5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            1   !       0   !       V   !    ]��     �   /   1   A      	         �   /   1   @    5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            2   !       1   !       V   !    ]��     �   2   5   B      	         �   2   4   A    5�_�   �   �           �   4        ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   3   5   C    �   4   5   C    5�_�   �   �           �   4   	    ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   4   6   E      	         �   4   6   D    5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   2   4   F      	         �   2   4   E    5�_�   �   �           �   5   	    ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   4   6          A         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);5�_�   �   �           �   6       ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   5   7                end if5�_�   �   �           �   7        ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   6   7           5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��     �   /   0          	         5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                            "   	       )   	       V   	    ]��     �   !   "             loop_proc: process      variable i: integer := 0;      begin         for i in 0 to 10 loop            wait for 320 ns;   A         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);         end loop;      end process;5�_�   �   �   �       �   +        ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]��   * �   +   -   =                  �   +   -   <    5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]��   + �   +   -   =                  i=0;5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]��   , �   -   /   =               end if5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]�
     �   *   ,   =               if(i=8) then5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]�     �   *   ,   =               if(i.=8) then5�_�   �   �           �   ,        ����                                                                                                                                                                                                                                                                                                                            (          )          V       ]�     �   +   .   =    �   ,   -   =    5�_�   �   �           �   -   	    ����                                                                                                                                                                                                                                                                                                                            (          )          V       ]�     �   -   /   @      	         �   -   /   ?    5�_�   �   �           �   (   	    ����                                                                                                                                                                                                                                                                                                                            )   	       (   	       V   	    ]�     �   '   (          %         spi_mosi_tb <= inData_tb(7);   4         inData_tb   <= inData_tb(6 downto 0) & '0';5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�     �   '   (                   i:=i+1;5�_�   �   �           �   .   	    ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�!     �   .   0   =    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�"     �   /   1   >    �   /   0   >    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�#     �   .   /           5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�.     �   '   )   >               if(i/=8) then5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            (   	       (   	       V   	    ]�B     �   '   )   >               if(i/=7) then5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /          /          V       ]��     �   .   /                   i:=i+1;5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            /          /          V       ]��     �   '   )   =    �   (   )   =    5�_�   �   �           �   .   	    ����                                                                                                                                                                                                                                                                                                                            0          0          V       ]��     �   -   /   >    �   .   /   >    5�_�   �   �           �   .   	    ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��     �   -   /          %         spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   *   "    ����                                                                                                                                                                                                                                                                                                                            +          *   "       V   "    ]��     �   *   ,          4         inData_tb   <= inData_tb(6 downto 0) & '0';�   )   +          %         spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            +          *   "       V   "    ]��     �   +   -          
      else5�_�   �   �           �   -        ����                                                                                                                                                                                                                                                                                                                            -   	       /   	       V   	    ]��   - �   <   >   ?      
        );�   ;   =   ?      !           clk          => clk_tb�   :   <   ?      '           ledsData     => ledsData_tb,�   9   ;   ?      '           inData       => inData_tb  ,�   8   :   ?      '           outData      => outData_tb ,�   7   9   ?      '           cs           => cs_tb      ,�   6   8   ?      '           spi_miso     => spi_miso_tb,�   5   7   ?      '    port map ( spi_mosi => spi_mosi_tb,�   4   6   ?         spi_inst: spi28b�   1   3   ?         end process;�   0   2   ?            end if;�   /   1   ?               end if;�   .   0   ?      F            inData_tb   <= std_logic_vector (unsigned(inData_tb) + 1);�   -   /   ?      (            spi_mosi_tb <= inData_tb(7);�   ,   .   ?                  i           := 0;�   +   -   ?               else�   *   ,   ?      7            inData_tb   <= inData_tb(6 downto 0) & '0';�   )   +   ?      (            spi_mosi_tb <= inData_tb(7);�   (   *   ?               if(i/=8) then�   '   )   ?               i:=i+1;�   &   (   ?      "      if rising_edge(clk_tb)  then�   %   '   ?         begin�   $   &   ?         �   #   %   ?         variable i :integer :=0;�   "   $   ?         spi_proc: process(clk_tb)�      !   ?         cs_tb    <= '0' after 1 ns;�          ?         rst_tb   <= '0';�         ?      &   clk_tb   <= not clk_tb after 20 ns;�         ?            �         ?      #    signal rst_tb      : STD_LOGIC;�         ?      *    signal clk_tb      : STD_LOGIC := '0';�         ?      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         ?      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         ?      7    signal outData_tb  : std_logic_vector (7 downto 0);�         ?      *    signal cs_tb       : std_logic := '1';�         ?      #    signal spi_miso_tb : STD_LOGIC;�         ?      #    signal spi_mosi_tb : STD_LOGIC;�         ?         end component;�         ?      
        );�         ?      %           clk      : in    STD_LOGIC�         ?      :           ledsData : out   std_logic_vector (3 downto 0);�         ?      :           inData   : in    std_logic_vector (7 downto 0);�         ?      :           outData  : out   std_logic_vector (7 downto 0);�         ?      &           cs       : in    std_logic;�   
      ?      &           spi_miso : out   STD_LOGIC;�   	      ?      &    port ( spi_mosi : in    STD_LOGIC;�      
   ?         component spi28b is�   ,   .                      i:=0;�   .   0          D            inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);�   -   /          (            spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   /   C    ����                                                                                                                                                                                                                                                                                                                            -   	       /   	       V   	    ]��   . �   .   0   ?      F            inData_tb   <= std_logic_vector (unsigned(inData_tb) + 1);5�_�   �   �           �   /   C    ����                                                                                                                                                                                                                                                                                                                            -   	       /   	       V   	    ]��   / �   .   0   ?      F            inData_tb   <= std_logic_vector (unsigned(inData_tb) + 2);5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                            -   	       /   	       V   	    ]�!     �         ?    �         ?    5�_�   �   �   �       �   %       ����                                                                                                                                                                                                                                                                                                                            .   	       0   	       V   	    ]�8     �   $   &   @    �   %   &   @    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            /   	       1   	       V   	    ]�:     �   %   '   A         variable i :integer :=0;5�_�   �   �           �   1   -    ����                                                                                                                                                                                                                                                                                                                            1   -       1   ?       v   ?    ]�C     �   0   2   A      F            inData_tb   <= std_logic_vector (unsigned(inData_tb) + 1);5�_�   �   �           �   1   /    ����                                                                                                                                                                                                                                                                                                                            1   -       1   ?       v   ?    ]�H     �   0   2   A      5            inData_tb   <= std_logic_vector (in + 1);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            1   -       1   ?       v   ?    ]�O     �   %   '   A         variable in :integer :=0;5�_�   �   �   �       �   %        ����                                                                                                                                                                                                                                                                                                                            &          %          V       ]�U     �   >   @   A      
        );�   =   ?   A      !           clk          => clk_tb�   <   >   A      '           ledsData     => ledsData_tb,�   ;   =   A      '           inData       => inData_tb  ,�   :   <   A      '           outData      => outData_tb ,�   9   ;   A      '           cs           => cs_tb      ,�   8   :   A      '           spi_miso     => spi_miso_tb,�   7   9   A      '    port map ( spi_mosi => spi_mosi_tb,�   6   8   A         spi_inst: spi28b�   3   5   A         end process;�   2   4   A            end if;�   1   3   A               end if;�   0   2   A      A            inData_tb   <= std_logic_vector (inData_integer + 1);�   /   1   A      (            spi_mosi_tb <= inData_tb(7);�   .   0   A                  i           := 0;�   -   /   A               else�   ,   .   A      7            inData_tb   <= inData_tb(6 downto 0) & '0';�   +   -   A      (            spi_mosi_tb <= inData_tb(7);�   *   ,   A               if(i/=8) then�   )   +   A               i:=i+1;�   (   *   A      "      if rising_edge(clk_tb)  then�   '   )   A         begin�   &   (   A         �   %   '   A      )   variable inData_integer :integer := 0;�   $   &   A      )   variable i :integer              := 0;�   #   %   A         spi_proc: process(clk_tb)�       "   A         cs_tb    <= '0' after 1 ns;�      !   A         rst_tb   <= '0';�          A      &   clk_tb   <= not clk_tb after 20 ns;�         A            �         A      #    signal rst_tb      : STD_LOGIC;�         A      *    signal clk_tb      : STD_LOGIC := '0';�         A      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         A      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         A      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         A      7    signal outData_tb  : std_logic_vector (7 downto 0);�         A      *    signal cs_tb       : std_logic := '1';�         A      #    signal spi_miso_tb : STD_LOGIC;�         A      #    signal spi_mosi_tb : STD_LOGIC;�         A         end component;�         A      
        );�         A      %           clk      : in    STD_LOGIC�         A      :           ledsData : out   std_logic_vector (3 downto 0);�         A      :           inData   : in    std_logic_vector (7 downto 0);�         A      :           outData  : out   std_logic_vector (7 downto 0);�         A      &           cs       : in    std_logic;�   
      A      &           spi_miso : out   STD_LOGIC;�   	      A      &    port ( spi_mosi : in    STD_LOGIC;�      
   A         component spi28b is�   $   &             variable i :integer :=0;�   %   '          (   variable inData_integer :integer :=0;5�_�   �   �   �       �   %       ����                                                                                                                                                                                                                                                                                                                            %           &           V        ]�]     �   $   &   A      )   variable i :integer              := 0;5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            %          &          V       ]�`   0 �   >   @   A      
        );�   =   ?   A      !           clk          => clk_tb�   <   >   A      '           ledsData     => ledsData_tb,�   ;   =   A      '           inData       => inData_tb  ,�   :   <   A      '           outData      => outData_tb ,�   9   ;   A      '           cs           => cs_tb      ,�   8   :   A      '           spi_miso     => spi_miso_tb,�   7   9   A      '    port map ( spi_mosi => spi_mosi_tb,�   6   8   A         spi_inst: spi28b�   3   5   A         end process;�   2   4   A            end if;�   1   3   A               end if;�   0   2   A      A            inData_tb   <= std_logic_vector (inData_integer + 1);�   /   1   A      (            spi_mosi_tb <= inData_tb(7);�   .   0   A                  i           := 0;�   -   /   A               else�   ,   .   A      7            inData_tb   <= inData_tb(6 downto 0) & '0';�   +   -   A      (            spi_mosi_tb <= inData_tb(7);�   *   ,   A               if(i/=8) then�   )   +   A               i:=i+1;�   (   *   A      "      if rising_edge(clk_tb)  then�   '   )   A         begin�   &   (   A         �   %   '   A      )   variable inData_integer :integer := 0;�   $   &   A      )   variable i              :integer := 0;�   #   %   A         spi_proc: process(clk_tb)�       "   A         cs_tb    <= '0' after 1 ns;�      !   A         rst_tb   <= '0';�          A      &   clk_tb   <= not clk_tb after 20 ns;�         A            �         A      #    signal rst_tb      : STD_LOGIC;�         A      *    signal clk_tb      : STD_LOGIC := '0';�         A      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         A      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         A      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         A      7    signal outData_tb  : std_logic_vector (7 downto 0);�         A      *    signal cs_tb       : std_logic := '1';�         A      #    signal spi_miso_tb : STD_LOGIC;�         A      #    signal spi_mosi_tb : STD_LOGIC;�         A         end component;�         A      
        );�         A      %           clk      : in    STD_LOGIC�         A      :           ledsData : out   std_logic_vector (3 downto 0);�         A      :           inData   : in    std_logic_vector (7 downto 0);�         A      :           outData  : out   std_logic_vector (7 downto 0);�         A      &           cs       : in    std_logic;�   
      A      &           spi_miso : out   STD_LOGIC;�   	      A      &    port ( spi_mosi : in    STD_LOGIC;�      
   A         component spi28b is�   $   &          6   variable i              :integer              := 0;�   %   '          )   variable inData_integer :integer := 0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            %          &          V       ]�i   1 �                E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";5�_�   �   �           �   0   -    ����                                                                                                                                                                                                                                                                                                                            $          %          V       ]�t     �   /   1   @      A            inData_tb   <= std_logic_vector (inData_integer + 1);5�_�   �   �           �   0   D    ����                                                                                                                                                                                                                                                                                                                            $          %          V       ]�{   2 �   /   1   @      J            inData_tb   <= std_logic_vector (unsigned(inData_integer + 1);5�_�   �   �           �   0   -    ����                                                                                                                                                                                                                                                                                                                            0   -       0   5       v   5    ]��     �   /   1   @      K            inData_tb   <= std_logic_vector (unsigned(inData_integer) + 1);5�_�   �   �           �   0   ;    ����                                                                                                                                                                                                                                                                                                                            0   -       0   5       v   5    ]��   3 �   /   1   @      B            inData_tb   <= std_logic_vector (inData_integer) + 1);5�_�   �   �           �   0   -    ����                                                                                                                                                                                                                                                                                                                            0   -       0   5       v   5    ]��     �   /   1   @      A            inData_tb   <= std_logic_vector (inData_integer + 1);5�_�   �   �           �   0   G    ����                                                                                                                                                                                                                                                                                                                            0   -       0   5       v   5    ]��     �   /   1   @      M            inData_tb   <= std_logic_vector (to_unsigned(inData_integer + 1);5�_�   �   �           �   0   G    ����                                                                                                                                                                                                                                                                                                                            0   -       0   5       v   5    ]��   5 �   /   1   @      N            inData_tb   <= std_logic_vector (to_unsigned(inData_integer) + 1);5�_�   �   �   �       �   0   O    ����                                                                                                                                                                                                                                                                                                                            0   H       0   \       v   \    ]��   6 �   /   1   @      d            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_integer'length) + 1);5�_�   �   �           �   /   '    ����                                                                                                                                                                                                                                                                                                                            0   -       0   .       v   .    ]��     �   /   1   A                  �   /   1   @    5�_�   �   �           �   0   ,    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   /   1   A      -            inData_integer:=inData_integer+1l5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   0   2   A      _            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length) + 1);5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   0   2   A      ^            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length)+ 1);5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   0   2   A      ]            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length) 1);5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   0   2   A      \            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length)1);5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��     �   0   2   A      [            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));5�_�   �   �           �   1   Y    ����                                                                                                                                                                                                                                                                                                                            1   -       1   .       v   .    ]��   8 �   0   2   A      Z            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length);5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /           /           V        ]��     �   .   /          (            spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            /           /           V        ]��     �   )   +   @    �   *   +   @    5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                            0           0           V        ]��     �   +   ,          (            spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            /           /           V        ]��   9 �   )   +          (            spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            0           .           V        ]�)>   : �   =   ?   @      
        );�   <   >   @      !           clk          => clk_tb�   ;   =   @      '           ledsData     => ledsData_tb,�   :   <   @      '           inData       => inData_tb  ,�   9   ;   @      '           outData      => outData_tb ,�   8   :   @      '           cs           => cs_tb      ,�   7   9   @      '           spi_miso     => spi_miso_tb,�   6   8   @      '    port map ( spi_mosi => spi_mosi_tb,�   5   7   @         spi_inst: spi28b�   2   4   @         end process;�   1   3   @            end if;�   0   2   @               end if;�   /   1   @      ^            inData_tb      <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   .   0   @      /            inData_integer := inData_integer+1;�   -   /   @                   i              := 0;�   ,   .   @               else�   +   -   @      7            inData_tb   <= inData_tb(6 downto 0) & '0';�   *   ,   @               if(i/=8) then�   )   +   @      %         spi_mosi_tb <= inData_tb(7);�   (   *   @               i:=i+1;�   '   )   @      "      if rising_edge(clk_tb)  then�   &   (   @         begin�   %   '   @         �   $   &   @      )   variable inData_integer :integer := 0;�   #   %   @      )   variable i              :integer := 0;�   "   $   @         spi_proc: process(clk_tb)�      !   @         cs_tb    <= '0' after 1 ns;�          @         rst_tb   <= '0';�         @      &   clk_tb   <= not clk_tb after 20 ns;�         @            �         @      #    signal rst_tb      : STD_LOGIC;�         @      *    signal clk_tb      : STD_LOGIC := '0';�         @      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         @      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         @      7    signal outData_tb  : std_logic_vector (7 downto 0);�         @      *    signal cs_tb       : std_logic := '1';�         @      #    signal spi_miso_tb : STD_LOGIC;�         @      #    signal spi_mosi_tb : STD_LOGIC;�         @         end component;�         @      
        );�         @      %           clk      : in    STD_LOGIC�         @      :           ledsData : out   std_logic_vector (3 downto 0);�         @      :           inData   : in    std_logic_vector (7 downto 0);�         @      :           outData  : out   std_logic_vector (7 downto 0);�         @      &           cs       : in    std_logic;�   
      @      &           spi_miso : out   STD_LOGIC;�   	      @      &    port ( spi_mosi : in    STD_LOGIC;�      
   @         component spi28b is�   -   /                      i           := 0;�   /   1          [            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   .   0          -            inData_integer:=inData_integer+1;5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                            0           .           V        ]�,c     �   6   9   @      '    port map ( spi_mosi => spi_mosi_tb,5�_�   �   �           �   9        ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�,m     �   =   ?          !           clk          => clk_tb�   <   >          '           ledsData     => ledsData_tb,�   ;   =          '           inData       => inData_tb  ,�   :   <          '           outData      => outData_tb ,�   9   ;          '           cs           => cs_tb      ,�   8   :          '           spi_miso     => spi_miso_tb,5�_�   �   �   �       �   8        ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�,u   ; �   >   @   A      
        );�   =   ?   A      "                clk      => clk_tb�   <   >   A      (                ledsData => ledsData_tb,�   ;   =   A      (                inData   => inData_tb  ,�   :   <   A      (                outData  => outData_tb ,�   9   ;   A      (                cs       => cs_tb      ,�   8   :   A      (                spi_miso => spi_miso_tb,�   7   9   A      (                spi_mosi => spi_mosi_tb,�   6   8   A          port map ( �   5   7   A         spi_inst: spi28b�   2   4   A         end process;�   1   3   A            end if;�   0   2   A               end if;�   /   1   A      ^            inData_tb      <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   .   0   A      /            inData_integer := inData_integer+1;�   -   /   A                   i              := 0;�   ,   .   A               else�   +   -   A      7            inData_tb   <= inData_tb(6 downto 0) & '0';�   *   ,   A               if(i/=8) then�   )   +   A      %         spi_mosi_tb <= inData_tb(7);�   (   *   A               i:=i+1;�   '   )   A      "      if rising_edge(clk_tb)  then�   &   (   A         begin�   %   '   A         �   $   &   A      )   variable inData_integer :integer := 0;�   #   %   A      )   variable i              :integer := 0;�   "   $   A         spi_proc: process(clk_tb)�      !   A         cs_tb    <= '0' after 1 ns;�          A         rst_tb   <= '0';�         A      &   clk_tb   <= not clk_tb after 20 ns;�         A            �         A      #    signal rst_tb      : STD_LOGIC;�         A      *    signal clk_tb      : STD_LOGIC := '0';�         A      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         A      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         A      7    signal outData_tb  : std_logic_vector (7 downto 0);�         A      *    signal cs_tb       : std_logic := '1';�         A      #    signal spi_miso_tb : STD_LOGIC;�         A      #    signal spi_mosi_tb : STD_LOGIC;�         A         end component;�         A      
        );�         A      %           clk      : in    STD_LOGIC�         A      :           ledsData : out   std_logic_vector (3 downto 0);�         A      :           inData   : in    std_logic_vector (7 downto 0);�         A      :           outData  : out   std_logic_vector (7 downto 0);�         A      &           cs       : in    std_logic;�   
      A      &           spi_miso : out   STD_LOGIC;�   	      A      &    port ( spi_mosi : in    STD_LOGIC;�      
   A         component spi28b is�   <   >          ,                ledsData     => ledsData_tb,�   ;   =          ,                inData       => inData_tb  ,�   7   9          (                spi_mosi => spi_mosi_tb,�   =   ?          &                clk          => clk_tb�   :   <          ,                outData      => outData_tb ,�   9   ;          ,                cs           => cs_tb      ,�   8   :          ,                spi_miso     => spi_miso_tb,5�_�   �   �           �   (   	    ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�1�   < �   '   )   A      "      if rising_edge(clk_tb)  then5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�1�   = �         A      *    signal clk_tb      : STD_LOGIC := '0';5�_�   �   �   �       �   *        ����                                                                                                                                                                                                                                                                                                                            ,           *           V        ]��     �   +   -          7            inData_tb   <= inData_tb(6 downto 0) & '0';�   )   +          %         spi_mosi_tb <= inData_tb(7);5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /          0          V       ]��#     �   .   1   A    �   /   0   A    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                            /          0          V       ]��(     �   /   1          ^            inData_tb      <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   .   0          /            inData_integer := inData_integer+1;5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            /          0          V       ]��5     �   $   &   C    �   %   &   C    5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            &          &          V       ]��7     �   %   '          )   variable inData_integer :integer := 0;5�_�   �   �           �   &   (    ����                                                                                                                                                                                                                                                                                                                            &          &          V       ]��9     �   %   '   D      *   variable outData_integer :integer := 0;5�_�   �   �           �   $        ����                                                                                                                                                                                                                                                                                                                            &   )       $   )       V   )    ]��?     �   A   C   D      
        );�   @   B   D      "                clk      => clk_tb�   ?   A   D      (                ledsData => ledsData_tb,�   >   @   D      (                inData   => inData_tb  ,�   =   ?   D      (                outData  => outData_tb ,�   <   >   D      (                cs       => cs_tb      ,�   ;   =   D      (                spi_miso => spi_miso_tb,�   :   <   D      (                spi_mosi => spi_mosi_tb,�   9   ;   D          port map ( �   8   :   D         spi_inst: spi28b�   5   7   D         end process;�   4   6   D            end if;�   3   5   D               end if;�   2   4   D      ^            inData_tb      <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   1   3   D      /            inData_integer := inData_integer+1;�   0   2   D      a            outData_tb      <= std_logic_vector (to_unsigned(outData_integer,outData_tb'length));�   /   1   D      1            outData_integer := outData_integer+1;�   .   0   D                   i              := 0;�   -   /   D               else�   ,   .   D      9            outData_tb   <= outData_tb(6 downto 0) & '0';�   +   -   D               if(i/=8) then�   *   ,   D      &         spi_mosi_tb <= outData_tb(7);�   )   +   D               i:=i+1;�   (   *   D      #      if falling_edge(clk_tb)  then�   '   )   D         begin�   &   (   D         �   %   '   D      ,   variable outData_integer :integer := 100;�   $   &   D      *   variable inData_integer :integer  := 0;�   #   %   D      *   variable i              :integer  := 0;�   "   $   D         spi_proc: process(clk_tb)�      !   D         cs_tb    <= '0' after 1 ns;�          D         rst_tb   <= '0';�         D      &   clk_tb   <= not clk_tb after 20 ns;�         D            �         D      #    signal rst_tb      : STD_LOGIC;�         D      *    signal clk_tb      : STD_LOGIC := '1';�         D      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         D      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         D      7    signal outData_tb  : std_logic_vector (7 downto 0);�         D      *    signal cs_tb       : std_logic := '1';�         D      #    signal spi_miso_tb : STD_LOGIC;�         D      #    signal spi_mosi_tb : STD_LOGIC;�         D         end component;�         D      
        );�         D      %           clk      : in    STD_LOGIC�         D      :           ledsData : out   std_logic_vector (3 downto 0);�         D      :           inData   : in    std_logic_vector (7 downto 0);�         D      :           outData  : out   std_logic_vector (7 downto 0);�         D      &           cs       : in    std_logic;�   
      D      &           spi_miso : out   STD_LOGIC;�   	      D      &    port ( spi_mosi : in    STD_LOGIC;�      
   D         component spi28b is�   #   %          )   variable i              :integer := 0;�   %   '          ,   variable outData_integer :integer := 100;�   $   &          )   variable inData_integer :integer := 0;5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            &          &          V       ]�ɬ     �   %   '          ,   variable outData_integer :integer := 100;5�_�   �              �   +        ����                                                                                                                                                                                                                                                                                                                            +          -          V       ]�ɳ     �   ,   .          9            outData_tb   <= outData_tb(6 downto 0) & '0';�   *   ,          &         spi_mosi_tb <= outData_tb(7);5�_�   �                0        ����                                                                                                                                                                                                                                                                                                                            0          1          V       ]�ɸ   > �   0   2          a            outData_tb      <= std_logic_vector (to_unsigned(outData_integer,outData_tb'length));�   /   1          1            outData_integer := outData_integer+1;5�_�                '        ����                                                                                                                                                                                                                                                                                                                            0          1          V       ]��     �   &   (   D    �   '   (   D    5�_�                 '       ����                                                                                                                                                                                                                                                                                                                            1          2          V       ]��     �   &   (   E      7    signal outData_tb  : std_logic_vector (7 downto 0);5�_�                 '       ����                                                                                                                                                                                                                                                                                                                            1          2          V       ]��      �   &   (   E      6    ignal outData_tb  : std_logic_vector (7 downto 0);5�_�                 '        ����                                                                                                                                                                                                                                                                                                                            '   
       '   
       V   
    ]��#   @ �   &   (          6   signal outData_tb  : std_logic_vector (7 downto 0);5�_�                 '        ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��/     �   &   '          7   signal mosiData_tb  : std_logic_vector (7 downto 0);5�_�    	                    ����                                                                                                                                                                                                                                                                                                                            '          '          V       ]��2     �         D    �         D    5�_�    
          	          ����                                                                                                                                                                                                                                                                                                                            (          (          V       ]��3     �         E    5�_�  	            
          ����                                                                                                                                                                                                                                                                                                                            )          )          V       ]��5   B �                7   signal mosiData_tb  : std_logic_vector (7 downto 0);5�_�  
                7    ����                                                                                                                                                                                                                                                                                                                            )          )          V       ]�ʀ   C �         F      8    signal mosiData_tb  : std_logic_vector (7 downto 0);5�_�                 1        ����                                                                                                                                                                                                                                                                                                                            1          5          V       ^��   D �   C   E   F      
        );�   B   D   F      "                clk      => clk_tb�   A   C   F      (                ledsData => ledsData_tb,�   @   B   F      (                inData   => inData_tb  ,�   ?   A   F      (                outData  => outData_tb ,�   >   @   F      (                cs       => cs_tb      ,�   =   ?   F      (                spi_miso => spi_miso_tb,�   <   >   F      (                spi_mosi => spi_mosi_tb,�   ;   =   F          port map ( �   :   <   F         spi_inst: spi28b�   7   9   F         end process;�   6   8   F            end if;�   5   7   F               end if;�   4   6   F      `            inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   3   5   F      1            inData_integer   := inData_integer+1;�   2   4   F      d            mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   1   3   F      3            mosiData_integer := mosiData_integer+1;�   0   2   F      "            i                := 0;�   /   1   F               else�   .   0   F      ;            mosiData_tb   <= mosiData_tb(6 downto 0) & '0';�   -   /   F               if(i/=8) then�   ,   .   F      '         spi_mosi_tb <= mosiData_tb(7);�   +   -   F               i:=i+1;�   *   ,   F      #      if falling_edge(clk_tb)  then�   )   +   F         begin�   (   *   F         �   '   )   F      -   variable mosiData_integer :integer := 100;�   &   (   F      *   variable inData_integer :integer  := 0;�   %   '   F      *   variable i              :integer  := 0;�   $   &   F         spi_proc: process(clk_tb)�   !   #   F         cs_tb    <= '0' after 1 ns;�       "   F         rst_tb   <= '0';�      !   F      &   clk_tb   <= not clk_tb after 20 ns;�         F            �         F      D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";�         F      #    signal rst_tb      : STD_LOGIC;�         F      *    signal clk_tb      : STD_LOGIC := '1';�         F      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         F      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         F      7    signal outData_tb  : std_logic_vector (7 downto 0);�         F      *    signal cs_tb       : std_logic := '1';�         F      #    signal spi_miso_tb : STD_LOGIC;�         F      #    signal spi_mosi_tb : STD_LOGIC;�         F         end component;�         F      
        );�         F      %           clk      : in    STD_LOGIC�         F      :           ledsData : out   std_logic_vector (3 downto 0);�         F      :           inData   : in    std_logic_vector (7 downto 0);�         F      :           outData  : out   std_logic_vector (7 downto 0);�         F      &           cs       : in    std_logic;�   
      F      &           spi_miso : out   STD_LOGIC;�   	      F      &    port ( spi_mosi : in    STD_LOGIC;�      
   F         component spi28b is�   0   2                       i              := 0;�   4   6          ^            inData_tb      <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   3   5          /            inData_integer := inData_integer+1;�   2   4          d            mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   1   3          3            mosiData_integer := mosiData_integer+1;5�_�                 &        ����                                                                                                                                                                                                                                                                                                                            &           (           V        ^�#     �   C   E   F      
        );�   B   D   F      "                clk      => clk_tb�   A   C   F      (                ledsData => ledsData_tb,�   @   B   F      (                inData   => inData_tb  ,�   ?   A   F      (                outData  => outData_tb ,�   >   @   F      (                cs       => cs_tb      ,�   =   ?   F      (                spi_miso => spi_miso_tb,�   <   >   F      (                spi_mosi => spi_mosi_tb,�   ;   =   F          port map ( �   :   <   F         spi_inst: spi28b�   7   9   F         end process;�   6   8   F            end if;�   5   7   F               end if;�   4   6   F      `            inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   3   5   F      1            inData_integer   := inData_integer+1;�   2   4   F      d            mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   1   3   F      3            mosiData_integer := mosiData_integer+1;�   0   2   F      "            i                := 0;�   /   1   F               else�   .   0   F      ;            mosiData_tb   <= mosiData_tb(6 downto 0) & '0';�   -   /   F               if(i/=8) then�   ,   .   F      '         spi_mosi_tb <= mosiData_tb(7);�   +   -   F               i:=i+1;�   *   ,   F      #      if falling_edge(clk_tb)  then�   )   +   F         begin�   (   *   F         �   '   )   F      -   variable mosiData_integer :integer := 100;�   &   (   F      +   variable inData_integer :integer   := 0;�   %   '   F      +   variable i              :integer   := 0;�   $   &   F         spi_proc: process(clk_tb)�   !   #   F         cs_tb    <= '0' after 1 ns;�       "   F         rst_tb   <= '0';�      !   F      &   clk_tb   <= not clk_tb after 20 ns;�         F            �         F      D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";�         F      #    signal rst_tb      : STD_LOGIC;�         F      *    signal clk_tb      : STD_LOGIC := '1';�         F      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         F      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         F      7    signal outData_tb  : std_logic_vector (7 downto 0);�         F      *    signal cs_tb       : std_logic := '1';�         F      #    signal spi_miso_tb : STD_LOGIC;�         F      #    signal spi_mosi_tb : STD_LOGIC;�         F         end component;�         F      
        );�         F      %           clk      : in    STD_LOGIC�         F      :           ledsData : out   std_logic_vector (3 downto 0);�         F      :           inData   : in    std_logic_vector (7 downto 0);�         F      :           outData  : out   std_logic_vector (7 downto 0);�         F      &           cs       : in    std_logic;�   
      F      &           spi_miso : out   STD_LOGIC;�   	      F      &    port ( spi_mosi : in    STD_LOGIC;�      
   F         component spi28b is�   %   '          *   variable i              :integer  := 0;�   &   (          *   variable inData_integer :integer  := 0;�   '   )          -   variable mosiData_integer :integer := 100;5�_�                 /        ����                                                                                                                                                                                                                                                                                                                            /           /           V        ^�)   E �   C   E   F      
        );�   B   D   F      "                clk      => clk_tb�   A   C   F      (                ledsData => ledsData_tb,�   @   B   F      (                inData   => inData_tb  ,�   ?   A   F      (                outData  => outData_tb ,�   >   @   F      (                cs       => cs_tb      ,�   =   ?   F      (                spi_miso => spi_miso_tb,�   <   >   F      (                spi_mosi => spi_mosi_tb,�   ;   =   F          port map ( �   :   <   F         spi_inst: spi28b�   7   9   F         end process;�   6   8   F            end if;�   5   7   F               end if;�   4   6   F      `            inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   3   5   F      1            inData_integer   := inData_integer+1;�   2   4   F      d            mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   1   3   F      3            mosiData_integer := mosiData_integer+1;�   0   2   F      "            i                := 0;�   /   1   F               else�   .   0   F      9            mosiData_tb <= mosiData_tb(6 downto 0) & '0';�   -   /   F               if(i/=8) then�   ,   .   F      '         spi_mosi_tb <= mosiData_tb(7);�   +   -   F               i:=i+1;�   *   ,   F      #      if falling_edge(clk_tb)  then�   )   +   F         begin�   (   *   F         �   '   )   F      -   variable mosiData_integer :integer := 100;�   &   (   F      +   variable inData_integer :integer   := 0;�   %   '   F      +   variable i              :integer   := 0;�   $   &   F         spi_proc: process(clk_tb)�   !   #   F         cs_tb    <= '0' after 1 ns;�       "   F         rst_tb   <= '0';�      !   F      &   clk_tb   <= not clk_tb after 20 ns;�         F            �         F      D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";�         F      #    signal rst_tb      : STD_LOGIC;�         F      *    signal clk_tb      : STD_LOGIC := '1';�         F      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         F      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         F      7    signal outData_tb  : std_logic_vector (7 downto 0);�         F      *    signal cs_tb       : std_logic := '1';�         F      #    signal spi_miso_tb : STD_LOGIC;�         F      #    signal spi_mosi_tb : STD_LOGIC;�         F         end component;�         F      
        );�         F      %           clk      : in    STD_LOGIC�         F      :           ledsData : out   std_logic_vector (3 downto 0);�         F      :           inData   : in    std_logic_vector (7 downto 0);�         F      :           outData  : out   std_logic_vector (7 downto 0);�         F      &           cs       : in    std_logic;�   
      F      &           spi_miso : out   STD_LOGIC;�   	      F      &    port ( spi_mosi : in    STD_LOGIC;�      
   F         component spi28b is�   .   0          ;            mosiData_tb   <= mosiData_tb(6 downto 0) & '0';5�_�                 A       ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^��     �   @   B   F      (                inData   => inData_tb  ,�   A   B   F    5�_�                 A   &    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^��   F �   @   B   F      2                inData   => outData_tbinData_tb  ,5�_�                 A   '    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�    G �   @   B   F      5                inData   => outData_tb;--inData_tb  ,5�_�                 A   &    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�/     �   @   B   F      7                inData   => outData_tb;  --inData_tb  ,5�_�                 A   &    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�0     �   @   B   F      8                inData   => outData_tb ;  --inData_tb  ,5�_�                 A   &    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�1     �   @   B   F      8                inData   => outData_tbl;  --inData_tb  ,5�_�                 A   &    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�3     �   @   B   F      8                inData   => outData_tb,;  --inData_tb  ,5�_�                 A   '    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�4     �   @   B   F      9                inData   => outData_tb ,;  --inData_tb  ,5�_�                 A   '    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�4     �   @   B   F      8                inData   => outData_tb ;  --inData_tb  ,5�_�                 A   '    ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�5   J �   @   B   F      7                inData   => outData_tb   --inData_tb  ,5�_�                       ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^��     �         F    �         F    5�_�                        ����                                                                                                                                                                                                                                                                                                                            A          A   %       v   %    ^��     �         G      #    signal rst_tb      : STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                            A          A   %       v   %    ^��     �         G          signal ii      : STD_LOGIC;5�_�                        ����                                                                                                                                                                                                                                                                                                                            A          A   %       v   %    ^��     �         G          signal ii      : integar;5�_�                         ����                                                                                                                                                                                                                                                                                                                            A          A   %       v   %    ^��     �         G          signal ii      : integer;5�_�    !              :        ����                                                                                                                                                                                                                                                                                                                            A          A   %       v   %    ^��     �   9   ;   G       5�_�     "          !   '        ����                                                                                                                                                                                                                                                                                                                            '          8          V       ^�     �   &   9   G      +   variable i              :integer   := 0;   +   variable inData_integer :integer   := 0;   -   variable mosiData_integer :integer := 100;            begin   #      if falling_edge(clk_tb)  then            i:=i+1;   '         spi_mosi_tb <= mosiData_tb(7);            if(i/=8) then   9            mosiData_tb <= mosiData_tb(6 downto 0) & '0';            else   "            i                := 0;   3            mosiData_integer := mosiData_integer+1;   d            mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));   1            inData_integer   := inData_integer+1;   `            inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));            end if;         end if;5�_�  !  #          "   :       ����                                                                                                                                                                                                                                                                                                                            '          8          V       ^�     �   9   ;   G        ii:=i5�_�  "  $          #   :        ����                                                                                                                                                                                                                                                                                                                            :          :          V       ^�
     �   9   :             ii:=i5�_�  #  %          $   9        ����                                                                                                                                                                                                                                                                                                                            :          :          V       ^�     �   8   :   F    �   9   :   F    5�_�  $  &          %   9       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^�   K �   8   :   G         ii:=i5�_�  %  '          &   9       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^�     �   8   :   G            ii:=i5�_�  &  (          '   9       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^��   L �   8   :   G            ii<=i5�_�  '  )          (      '    ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^�s   M �         G      *    signal clk_tb      : STD_LOGIC := '1';5�_�  (  *          )      '    ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^��   N �         G      *    signal clk_tb      : STD_LOGIC := '0';5�_�  )  +          *   #       ����                                                                                                                                                                                                                                                                                                                            ;          ;          V       ^��   O �   "   $   G         cs_tb    <= '0' after 1 ns;5�_�  *  ,          +   #       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�     �   "   $   G         cs_tb    <= '0' after 5 ns;�   #   $   G    5�_�  +  -          ,   #   %    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�     �   "   %   G      4   cs_tb    <= not clk_tb after 20 ns'0' after 5 ns;5�_�  ,  .          -   #       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�     �   "   $   H      %   cs_tb    <= not clk_tb after 20 ns5�_�  -  /          .   #       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�   P �   "   $   H      $   cs_tb    <= not cs_tb after 20 ns5�_�  .  0          /   #   %    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�&   R �   "   $   H      %   cs_tb    <= not cs_tb after 160 ns5�_�  /  1          0   #        ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�e     �   "   $   H      &   cs_tb    <= not cs_tb after 160 ns;5�_�  0  2          1   #   !    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�f     �   "   $   H      &   cs_tb    <= not cs_tb after 150 ns;5�_�  1  3          2   #   !    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^�i   S �   "   $   H      &   cs_tb    <= not cs_tb after 159 ns;5�_�  2  4          3   #       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��   T �   "   $   H      &   cs_tb    <= not cs_tb after 155 ns;5�_�  3  5          4      6    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �         H      7    signal outData_tb  : std_logic_vector (7 downto 0);5�_�  4  6          5      C    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �         H      E    signal outData_tb  : std_logic_vector (7 downto 0) := '01010101';5�_�  5  7          6      :    ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��   U �         H      E    signal outData_tb  : std_logic_vector (7 downto 0) := '01010101";5�_�  6  8          7   *        ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   *   -   I            �   *   ,   H    5�_�  7  9          8   ,        ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   ,   .   J    �   ,   -   J    5�_�  8  :          9   ,        ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   +   ,           5�_�  9  ;          :   ,       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   +   -   J            cs_tb <= '1'5�_�  :  <          ;   ,       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   +   -   J            cs_tb <= '0'5�_�  ;  =          <   ,       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��     �   +   -   J            cs_tb <= '0' after 100ns5�_�  <  >          =   ,       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��   V �   +   -   J            cs_tb <= '0' after 100 ns5�_�  =  ?          >   +       ����                                                                                                                                                                                                                                                                                                                            !          !   $       v   $    ^��   W �   *   ,   J            cs_tb <= '1'5�_�  >  @          ?   +        ����                                                                                                                                                                                                                                                                                                                            +          -          V       ^��     �   *   +                cs_tb <= '1';          cs_tb <= '0' after 100 ns;         5�_�  ?  A          @   ,       ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^��     �   +   /   G    �   ,   -   G    5�_�  @  B          A   +       ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^��     �   +   -   J    5�_�  A  C          B   *   	    ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^��     �   *   ,   K    5�_�  B  D          C   -        ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^��     �   ,   -           5�_�  C  E          D   -        ����                                                                                                                                                                                                                                                                                                                            -          .          V       ^��   X �   -   /                 cs_tb <= '0' after 100 ns;�   ,   .                cs_tb <= '1';5�_�  D  F          E   -        ����                                                                                                                                                                                                                                                                                                                            -           .           V        ^�     �   ,   -                   cs_tb <= '1';   #         cs_tb <= '0' after 100 ns;5�_�  E  G          F   &        ����                                                                                                                                                                                                                                                                                                                            -           -           V        ^�	     �   %   (   I    �   &   '   I    5�_�  F  H          G   &        ����                                                                                                                                                                                                                                                                                                                            &          '          V       ^�!     �   %   &                   cs_tb <= '1';   #         cs_tb <= '0' after 100 ns;5�_�  G  I          H   -        ����                                                                                                                                                                                                                                                                                                                            &          &          V       ^�:     �   ,   -                5�_�  H  J          I   -   	    ����                                                                                                                                                                                                                                                                                                                            &          &          V       ^�;     �   -   /   I                  �   -   /   H    5�_�  I  K          J   /        ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�N     �   .   :   I                  i:=i+1;   *            spi_mosi_tb <= mosiData_tb(7);               if(i/=8) then   <               mosiData_tb <= mosiData_tb(6 downto 0) & '0';               else   %               i                := 0;   6               mosiData_integer := mosiData_integer+1;   g               mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));   4               inData_integer   := inData_integer+1;   c               inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));               end if;5�_�  J  L          K   9       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�Q   Y �   9   <   J                     �   9   ;   I    5�_�  K  M          L   <       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�]     �   ;   =   K    �   <   =   K    5�_�  L  N          M   <   	    ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�_   Z �   ;   =                   end if;5�_�  M  O          N   <       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^��     �   ;   =   L    �   <   =   L    5�_�  N  P          O   <       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^��     �   ;   =   M      j                  mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));5�_�  O  Q          P   <       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^��     �   ;   =   M      i                 mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));5�_�  P  R          Q   <       ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^��   [ �   ;   =   M      h                mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));5�_�  Q  S          R   #        ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�s     �   "   $   M      &   cs_tb    <= not cs_tb after 317 ns;5�_�  R  T          S      '    ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^��   \ �         M      *    signal clk_tb      : STD_LOGIC := '1';5�_�  S  V          T   ,   
    ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�;     �   ,   .   N      	         �   ,   .   M    5�_�  T  W  U      V   -   	    ����                                                                                                                                                                                                                                                                                                                            0          :          V       ^�U     �   ,   -                   wait for 1005�_�  V  X          W   &        ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�W     �   %   )   M       5�_�  W  Y          X   '        ����                                                                                                                                                                                                                                                                                                                            1          ;          V       ^�X     �   &   +   O       5�_�  X  Z          Y   +        ����                                                                                                                                                                                                                                                                                                                            4          >          V       ^�~     �   *   ,   R    �   +   ,   R    5�_�  Y  [          Z   +       ����                                                                                                                                                                                                                                                                                                                            5          ?          V       ^�     �   +   -   T            �   +   -   S    5�_�  Z  \          [   #        ����                                                                                                                                                                                                                                                                                                                            6          @          V       ^��   ] �   "   $   T      &   cs_tb    <= not cs_tb after 320 ns;5�_�  [  ]          \   '       ����                                                                                                                                                                                                                                                                                                                            6          @          V       ^��   ^ �   '   )   U            �   '   )   T    5�_�  \  ^          ]   *       ����                                                                                                                                                                                                                                                                                                                            7          A          V       ^��     �   )   +   U            wait for 100ns;5�_�  ]  _          ^   ,       ����                                                                                                                                                                                                                                                                                                                            7          A          V       ^��   _ �   +   -   U            wait for 100ns;5�_�  ^  `          _   -       ����                                                                                                                                                                                                                                                                                                                            7          A          V       ^��   ` �   ,   .   U         end process5�_�  _  a          `   ,       ����                                                                                                                                                                                                                                                                                                                            7          A          V       ^��     �   ,   /   V            �   ,   .   U    5�_�  `  b          a   -       ����                                                                                                                                                                                                                                                                                                                            9          C          V       ^�(     �   ,   .   W            for k in 0 to 8 loop5�_�  a  c          b   .       ����                                                                                                                                                                                                                                                                                                                            9          C          V       ^�/     �   -   /   W               end loop5�_�  b  d          c   -       ����                                                                                                                                                                                                                                                                                                                            9          C          V       ^�2     �   -   /   X      	         �   -   /   W    5�_�  c  e          d   .   	    ����                                                                                                                                                                                                                                                                                                                            :          D          V       ^�5     �   -   /   X      
         j5�_�  d  f          e   .   	    ����                                                                                                                                                                                                                                                                                                                            :          D          V       ^�9     �   -   0   X      	         5�_�  e  g          f   .   	    ����                                                                                                                                                                                                                                                                                                                            ;          E          V       ^�N     �   -   /   Y    5�_�  f  h          g   .        ����                                                                                                                                                                                                                                                                                                                            <          F          V       ^�R     �   -   /   [      	         �   -   /   Z    5�_�  g  i          h   .        ����                                                                                                                                                                                                                                                                                                                            .   	       .   	       V   	    ^�Y     �   -   /   Z    �   .   /   Z    �   -   .          
         h5�_�  h  j          i   1        ����                                                                                                                                                                                                                                                                                                                            .           .          V   	    ^�]     �   0   2   [    5�_�  i  k          j   1        ����                                                                                                                                                                                                                                                                                                                            .           .          V   	    ^�`     �   0   2   \    �   1   2   \    5�_�  j  l          k   /        ����                                                                                                                                                                                                                                                                                                                            .           .          V   	    ^�b     �   .   /           5�_�  k  m          l   /   	    ����                                                                                                                                                                                                                                                                                                                            .           .          V   	    ^�c     �   .   0                   clk_tb <= not clk_tb;5�_�  l  n          m   .        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�e     �   -   1   \            wait for 100 ns;         clk_tb <= not clk_tb;         wait for 100 ns;5�_�  m  o          n   0   	    ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�o     �   /   0                   wait for 100 ns;5�_�  n  p          o   0        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�o     �   /   0           5�_�  o  q          p   0        ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�p     �   /   0           5�_�  p  r          q   0   	    ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�s     �   /   1                   end loop clk_loop5�_�  q  s          r   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�w     �   ,   .   Y      #      clk_loop:for k in 0 to 8 loop5�_�  r  t          s   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^�     �   ,   .   Y      %      clk_loop:for k in 0 to 158 loop5�_�  s  u          t   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   ,   .   Y      %      clk_loop:for k in 0 to 108 loop5�_�  t  v          u   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   ,   .   Y      %      clk_loop:for k in 0 to 168 loop5�_�  u  w          v   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   ,   .   Y      %      clk_loop:for k in 0 to 168 loop5�_�  v  x          w   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   ,   .   Y      %      clk_loop:for k in 0 to 158 loop5�_�  w  y          x   -       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   ,   .   Y      %      clk_loop:for k in 0 to 168 loop5�_�  x  z          y   )       ����                                                                                                                                                                                                                                                                                                                            .          0          V       ^��     �   (   *   Y    �   )   *   Y    5�_�  y  {          z   )       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   (   *   Z            cs_tb <= '1';5�_�  z  |          {   )       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   (   *   Z            cl_tb <= '1';5�_�  {  }          |   )       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   (   *   Z            clk_tb <= '1';5�_�  |  ~          }   2       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   Z    �   2   3   Z    5�_�  }            ~   2       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   [    5�_�  ~  �             2        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   \    �   2   3   \    5�_�    �          �   2       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   ]               wait for 100 ns;5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   ]              wait for 100 ns;5�_�  �  �          �   2       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   1   3   ]             wait for 100 ns;5�_�  �  �          �   3        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   2   4   ]       5�_�  �  �          �   3        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   2   3           5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   3   5   \    5�_�  �  �          �   4        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   3   5   ]    5�_�  �  �          �   4        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   3   5   ^    �   4   5   ^    5�_�  �  �          �   4       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   3   5   _            wait for 100 ns;5�_�  �  �          �   5        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��     �   4   5           5�_�  �  �          �   5        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��   a �   4   5           5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��   b �   0   2   ]            end loop clk_loop5�_�  �  �          �   !        ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��   c �       "   ]      &   clk_tb   <= not clk_tb after 20 ns;5�_�  �  �          �   .       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^�6   d �   -   /   ]      $      clk_loop:for k in 0 to 16 loop5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                            /          1          V       ^��   e �   (   *   ]            clk_tb <= '0';5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      "                clk      => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      &                spi_clk      => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      %                spi_clk     => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      $                spi_clk    => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      #                spi_clk   => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      "                spi_clk  => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]      !                spi_clk => clk_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ]    �   Z   [   ]    5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^      "                spi_clk  => clk_tb5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^      !                pi_clk  => clk_tb5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^      "                sys_clk  => clk_tb5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^      !                sys_clk  => lk_tb5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^                       sys_clk  => k_tb5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^                      sys_clk  => _tb5�_�  �  �          �   [        ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Z   \   ^      "                sys_clk  => sys_tb5�_�  �  �          �   Z       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ^      "                spi_clk  => clk_tb5�_�  �  �          �   Z   &    ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   Y   [   ^      &                spi_clk  => spi_clk_tb5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   6   8   ^         spi_proc: process(clk_tb)5�_�  �  �          �   1       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   0   2   ^            end loop clk_loop;5�_�  �  �          �   0       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   /   1   ^               clk_tb <= not clk_tb;5�_�  �  �          �   0   	    ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   /   1   ^      "         clk_tb <= not spi_clk_tb;5�_�  �  �          �   .       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   -   /   ^      $      clk_loop:for k in 0 to 15 loop5�_�  �  �          �   )       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   (   *   ^            clk_tb <= '1';5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �       "   ^      (--   clk_tb   <= not clk_tb after 20 ns;5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �       "   ^      ,--   clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �         ^      *    signal clk_tb      : STD_LOGIC := '0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �         ^      %           clk      : in    STD_LOGIC5�_�  �  �          �   =       ����                                                                                                                                                                                                                                                                                                                                                             ^A�     �   <   >   ^      &         if falling_edge(clk_tb)  then5�_�  �  �          �   )        ����                                                                                                                                                                                                                                                                                                                            )   
       *   
       V   
    ^A�   f �   [   ]   ^      
        );�   Z   \   ^      &                sys_clk  => sys_clk_tb�   Y   [   ^      '                spi_clk  => spi_clk_tb,�   X   Z   ^      (                ledsData => ledsData_tb,�   W   Y   ^      7                inData   => outData_tb , --inData_tb  ,�   V   X   ^      (                outData  => outData_tb ,�   U   W   ^      (                cs       => cs_tb      ,�   T   V   ^      (                spi_miso => spi_miso_tb,�   S   U   ^      (                spi_mosi => spi_mosi_tb,�   R   T   ^          port map ( �   Q   S   ^         spi_inst: spi28b�   O   Q   ^         end process;�   N   P   ^            ii<=i;�   M   O   ^               end if;�   L   N   ^                  end if;�   K   M   ^      g               mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   J   L   ^                     i:=0;�   I   K   ^                  else �   H   J   ^                     end if;�   G   I   ^      f                  inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   F   H   ^      7                  inData_integer   := inData_integer+1;�   E   G   ^      j                  mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   D   F   ^      9                  mosiData_integer := mosiData_integer+1;�   C   E   ^      (                  i                := 0;�   B   D   ^                     else�   A   C   ^      ?                  mosiData_tb <= mosiData_tb(6 downto 0) & '0';�   @   B   ^                     if(i/=8) then�   ?   A   ^      -               spi_mosi_tb <= mosiData_tb(7);�   >   @   ^                     i:=i+1;�   =   ?   ^                  if cs_tb = '0' then�   <   >   ^      *         if falling_edge(spi_clk_tb)  then�   ;   =   ^            begin�   9   ;   ^      0      variable mosiData_integer :integer := 100;�   8   :   ^      .      variable inData_integer :integer   := 0;�   7   9   ^      .      variable i              :integer   := 0;�   6   8   ^          spi_proc: process(spi_clk_tb)�   4   6   ^         end process;�   3   5   ^            wait for 1000 ns;�   2   4   ^            cs_tb <= '1';�   1   3   ^            wait for 100 ns;�   0   2   ^            end loop spi_clk_loop;�   /   1   ^      &         spi_clk_tb <= not spi_clk_tb;�   .   0   ^               wait for 100 ns;�   -   /   ^      (      spi_clk_loop:for k in 0 to 15 loop�   ,   .   ^            wait for 100 ns;�   +   -   ^            cs_tb<='0';�   *   ,   ^            wait for 100 ns;�   )   +   ^            cs_tb      <= '1';�   (   *   ^            spi_clk_tb <= '1';�   '   )   ^         begin�   &   (   ^         cs_proc: process is�   #   %   ^                      --'0' after 5 ns;�   "   $   ^      (--   cs_tb    <= not cs_tb after 320 ns;�   !   #   ^         rst_tb   <= '0';�       "   ^      0--   spi_clk_tb   <= not spi_clk_tb after 20 ns;�          ^            �         ^      D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";�         ^      !    signal ii          : integer;�         ^      #    signal rst_tb      : STD_LOGIC;�         ^      .    signal spi_clk_tb      : STD_LOGIC := '0';�         ^      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         ^      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         ^      E    signal outData_tb  : std_logic_vector (7 downto 0) := "01010101";�         ^      *    signal cs_tb       : std_logic := '1';�         ^      #    signal spi_miso_tb : STD_LOGIC;�         ^      #    signal spi_mosi_tb : STD_LOGIC;�         ^         end component;�         ^      
        );�         ^      )           spi_clk      : in    STD_LOGIC�         ^      :           ledsData : out   std_logic_vector (3 downto 0);�         ^      :           inData   : in    std_logic_vector (7 downto 0);�         ^      :           outData  : out   std_logic_vector (7 downto 0);�         ^      &           cs       : in    std_logic;�   
      ^      &           spi_miso : out   STD_LOGIC;�   	      ^      &    port ( spi_mosi : in    STD_LOGIC;�      
   ^         component spi28b is�   (   *                spi_clk_tb <= '1';�   )   +                cs_tb <= '1';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            )   
       *   
       V   
    ^B,     �         ^      .    signal spi_clk_tb      : STD_LOGIC := '0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            )   
       *   
       V   
    ^B-     �         ^    �         ^    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^B/     �         _      *    signal spi_clk_tb  : STD_LOGIC := '0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^B/     �         _      )    signal pi_clk_tb  : STD_LOGIC := '0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^B/     �         _      (    signal i_clk_tb  : STD_LOGIC := '0';5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^B0   g �         _      '    signal _clk_tb  : STD_LOGIC := '0';5�_�  �  �  �      �   T       ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^BD   i �   S   U   _          port map ( 5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^Bs     �         _      )           spi_clk      : in    STD_LOGIC5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^Bt     �         _    �         _    5�_�  �  �          �      %    ����                                                                                                                                                                                                                                                                                                                            +   
       ,   
       V   
    ^Bv     �         `      %           spi_clk  : in    STD_LOGIC5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            +   
       ,   
       V   
    ^Bx   j �         `      %           spi_clk  : in    STD_LOGIC5�_�  �  �          �      %    ����                                                                                                                                                                                                                                                                                                                            +   
       ,   
       V   
    ^B   k �         `      &           spi_clk  : in    STD_LOGIC,5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                            +   
       ,   
       V   
    ^B�   m �   T   V   `          port map (5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            +   
       ,   
       V   
    ^B�     �   
      `    �         `    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ,   
       -   
       V   
    ^B�     �         a      &           spi_miso : out   STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       ^B�     �         a      %           pi_miso : out   STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       ^B�     �         a      '           stop_data : out   STD_LOGIC;5�_�  �  �          �   Y       ����                                                                                                                                                                                                                                                                                                                                                v       ^Cp     �   X   Z   a    �   Y   Z   a    5�_�  �  �          �   Y       ����                                                                                                                                                                                                                                                                                                                                                v       ^Cr     �   X   Z   b      &           stop_data: out   STD_LOGIC;5�_�  �  �          �   Y       ����                                                                                                                                                                                                                                                                                                                                                v       ^Cw     �   X   Z   b      +                stop_data: out   STD_LOGIC;5�_�  �  �          �   Y   (    ����                                                                                                                                                                                                                                                                                                                                                v       ^C�     �   X   Z   b      ;                stop_data => stop_data_tb: out   STD_LOGIC;5�_�  �  �          �   Y   )    ����                                                                                                                                                                                                                                                                                                                            Y   )       Y   9       v   9    ^C�     �   X   Z   b      ;                stop_data => stop_data_tb: out   STD_LOGIC;5�_�  �  �          �   W        ����                                                                                                                                                                                                                                                                                                                            W   '       `   
       V   )    ^C�   n �   _   a   b      
        );�   ^   `   b      '                sys_clk   => sys_clk_tb�   ]   _   b      (                spi_clk   => spi_clk_tb,�   \   ^   b      )                ledsData  => ledsData_tb,�   [   ]   b      8                inData    => outData_tb , --inData_tb  ,�   Z   \   b      )                outData   => outData_tb ,�   Y   [   b      )                cs        => cs_tb      ,�   X   Z   b      *                stop_data => stop_data_tb;�   W   Y   b      )                spi_miso  => spi_miso_tb,�   V   X   b      )                spi_mosi  => spi_mosi_tb,�   U   W   b         port map (�   T   V   b         spi_inst: spi28b�   R   T   b         end process;�   Q   S   b            ii<=i;�   P   R   b               end if;�   O   Q   b                  end if;�   N   P   b      g               mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   M   O   b                     i:=0;�   L   N   b                  else �   K   M   b                     end if;�   J   L   b      f                  inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));�   I   K   b      7                  inData_integer   := inData_integer+1;�   H   J   b      j                  mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));�   G   I   b      9                  mosiData_integer := mosiData_integer+1;�   F   H   b      (                  i                := 0;�   E   G   b                     else�   D   F   b      ?                  mosiData_tb <= mosiData_tb(6 downto 0) & '0';�   C   E   b                     if(i/=8) then�   B   D   b      -               spi_mosi_tb <= mosiData_tb(7);�   A   C   b                     i:=i+1;�   @   B   b                  if cs_tb = '0' then�   ?   A   b      *         if falling_edge(spi_clk_tb)  then�   >   @   b            begin�   <   >   b      0      variable mosiData_integer :integer := 100;�   ;   =   b      .      variable inData_integer :integer   := 0;�   :   <   b      .      variable i              :integer   := 0;�   9   ;   b          spi_proc: process(spi_clk_tb)�   7   9   b         end process;�   6   8   b            wait for 1000 ns;�   5   7   b            cs_tb <= '1';�   4   6   b            wait for 100 ns;�   3   5   b            end loop spi_clk_loop;�   2   4   b      &         spi_clk_tb <= not spi_clk_tb;�   1   3   b               wait for 100 ns;�   0   2   b      (      spi_clk_loop:for k in 0 to 15 loop�   /   1   b            wait for 100 ns;�   .   0   b            cs_tb<='0';�   -   /   b            wait for 100 ns;�   ,   .   b            cs_tb      <= '1';�   +   -   b            spi_clk_tb <= '1';�   *   ,   b         begin�   )   +   b         cs_proc: process is�   &   (   b                      --'0' after 5 ns;�   %   '   b      (--   cs_tb    <= not cs_tb after 320 ns;�   $   &   b         rst_tb   <= '0';�   #   %   b      0--   spi_clk_tb   <= not spi_clk_tb after 20 ns;�   !   #   b            �       "   b      D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";�          b      !    signal ii          : integer;�         b      #    signal rst_tb      : STD_LOGIC;�         b      *    signal sys_clk_tb  : STD_LOGIC := '0';�         b      *    signal spi_clk_tb  : STD_LOGIC := '0';�         b      7    signal ledsData_tb : std_logic_vector (3 downto 0);�         b      E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";�         b      E    signal outData_tb  : std_logic_vector (7 downto 0) := "01010101";�         b      *    signal cs_tb       : std_logic := '1';�         b      #    signal spi_miso_tb : STD_LOGIC;�         b      #    signal spi_mosi_tb : STD_LOGIC;�         b         end component;�         b      
        );�         b      %           sys_clk  : in    STD_LOGIC�         b      &           spi_clk  : in    STD_LOGIC;�         b      :           ledsData : out   std_logic_vector (3 downto 0);�         b      :           inData   : in    std_logic_vector (7 downto 0);�         b      :           outData  : out   std_logic_vector (7 downto 0);�         b      &           cs       : in    std_logic;�         b      &           stop_data: out   STD_LOGIC;�   
      b      &           spi_miso : out   STD_LOGIC;�   	      b      &    port ( spi_mosi : in    STD_LOGIC;�      
   b         component spi28b is�   [   ]          7                inData   => outData_tb , --inData_tb  ,�   Z   \          (                outData  => outData_tb ,�   Y   [          (                cs       => cs_tb      ,�   \   ^          (                ledsData => ledsData_tb,�   V   X          (                spi_mosi => spi_mosi_tb,�   ]   _          '                spi_clk  => spi_clk_tb,�   ^   `          &                sys_clk  => sys_clk_tb�   X   Z          *                stop_data => stop_data_tb;�   W   Y          (                spi_miso => spi_miso_tb,5�_�  �  �          �   Y   )    ����                                                                                                                                                                                                                                                                                                                            W   '       `   
       V   )    ^C�   o �   X   Z   b      *                stop_data => stop_data_tb;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            W   '       `   
       V   )    ^C�     �         b    �         b    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            X   '       a   
       V   )    ^C�     �         c      #    signal spi_miso_tb : STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       ^C�   p �         c      "    signal pi_miso_tb : STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                       ^C�     �         c      #    signal spi_miso_tb : STD_LOGIC;�         c      #    signal spi_mosi_tb : STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                        ^C�   r �      !   c      E    signal outData_tb  : std_logic_vector (7 downto 0) := "01010101";   E    signal inData_tb   : std_logic_vector (7 downto 0) := "00000000";   7    signal ledsData_tb : std_logic_vector (3 downto 0);   *    signal spi_clk_tb  : STD_LOGIC := '0';   *    signal sys_clk_tb  : STD_LOGIC := '0';   #    signal rst_tb      : STD_LOGIC;   !    signal ii          : integer;�         c      *    signal cs_tb       : std_logic := '1';5�_�  �  �          �   %        ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      0--   spi_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �          �   %        ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      /-   spi_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �  �      �   %       ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      .   spi_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �          �   %       ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      .   sys_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �          �   %   (    ����                                                                                                                                                                                                                                                                                                                                                        ^J�   s �   $   &   c      .   sys_clk_tb   <= not sys_clk_tb after 20 ns;5�_�  �  �          �   %   (    ����                                                                                                                                                                                                                                                                                                                                                             ^W�     �   $   &   c      .   sys_clk_tb   <= not sys_clk_tb after 15 ns;5�_�  �  �          �   %   +    ����                                                                                                                                                                                                                                                                                                                                                             ^W�     �   $   &   c      1   sys_clk_tb   <= not sys_clk_tb after 10015 ns;5�_�  �  �          �   %   ,    ����                                                                                                                                                                                                                                                                                                                                                             ^W�     �   $   &   c      2   sys_clk_tb   <= not sys_clk_tb after 100 15 ns;5�_�  �  �          �   %   ,    ����                                                                                                                                                                                                                                                                                                                                                             ^W�     �   $   &   c      1   sys_clk_tb   <= not sys_clk_tb after 100 5 ns;5�_�  �  �          �   %   ,    ����                                                                                                                                                                                                                                                                                                                                                             ^W�   t �   $   &   c      0   sys_clk_tb   <= not sys_clk_tb after 100  ns;5�_�  �  �          �   %   /    ����                                                                                                                                                                                                                                                                                                                                                             ^X   u �   $   &   c      /   sys_clk_tb   <= not sys_clk_tb after 100 ns;5�_�  �  �          �   %   3    ����                                                                                                                                                                                                                                                                                                                                                             ^X�     �   $   &   c      7   sys_clk_tb   <= not sys_clk_tb after 100 ns; --19Mhz5�_�  �  �          �   %   3    ����                                                                                                                                                                                                                                                                                                                                                             ^X�   v �   $   &   c      7   sys_clk_tb   <= not sys_clk_tb after 100 ns; --19Mhz5�_�  �  �  �      �   V       ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   U   W   c         spi_inst: spi28b5�_�  �  �          �   V        ����                                                                                                                                                                                                                                                                                                                            V           a           V        ^0      �   U   e   W    �   V   W   W    �   U   V             stretcher: spi28b      port map (   )                spi_mosi  => spi_mosi_tb,   )                spi_miso  => spi_miso_tb,   *                stop_data => stop_data_tb,   )                cs        => cs_tb      ,   )                outData   => outData_tb ,   8                inData    => outData_tb , --inData_tb  ,   )                ledsData  => ledsData_tb,   (                spi_clk   => spi_clk_tb,   '                sys_clk   => sys_clk_tb   
        );5�_�  �  �          �   W       ����                                                                                                                                                                                                                                                                                                                            V           d          V        ^0     �   V   X   f          Port(  5�_�  �  �          �   W       ����                                                                                                                                                                                                                                                                                                                            V           d          V        ^0     �   V   X   f          port(  5�_�  �  �          �   X        ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^0     �   b   d          *           rst           : in  STD_LOGIC);�   a   c          )           clk           : in  STD_LOGIC;�   _   a          )           s_axis_tready : out STD_LOGIC;�   ^   `          )           s_axis_tlast  : in  STD_LOGIC;�   ]   _          )           s_axis_tvalid : in  STD_LOGIC;�   \   ^          =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   Z   \          )           m_axis_tready : in  STD_LOGIC;�   Y   [          )           m_axis_tlast  : out STD_LOGIC;�   X   Z          )           m_axis_tvalid : out STD_LOGIC;�   W   Y          =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �   d        ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^0     �   c   d          end stretcher;5�_�  �  �          �   V        ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^0     �   U   W   e      entity stretcher is5�_�  �  �          �   V        ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^0     �   U   W   e      stretcher is5�_�  �  �          �   V       ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^07     �   U   W   e      stretcher_inst:stretcher is5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            X          c          V       ^0e     �      
   e    5�_�  �  �          �   	        ����                                                                                                                                                                                                                                                                                                                            Y          d          V       ^0e     �   	      f    �   	   
   f    5�_�  �  �          �   
        ����                                                                                                                                                                                                                                                                                                                            h          s          V       ^0f     �   	      u      entity stretcher is5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            h          s          V       ^0m     �   
      u          Port(  5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            h          s          V       ^0u     �         v          �         u    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       ^0�     �         v         end component;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                      %          V       ^0�     �                end stretcher;      component spi28b is   &    port ( spi_mosi : in    STD_LOGIC;   &           spi_miso : out   STD_LOGIC;   &           stop_data: out   STD_LOGIC;   &           cs       : in    std_logic;   :           outData  : out   std_logic_vector (7 downto 0);   :           inData   : in    std_logic_vector (7 downto 0);   :           ledsData : out   std_logic_vector (3 downto 0);   &           spi_clk  : in    STD_LOGIC;   %           sys_clk  : in    STD_LOGIC   
        );      end component;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                V       ^0�     �      #   i    �         i    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                      "                 ^0�     �      #   r      )           m_axis_tvalid : out STD_LOGIC;   )           m_axis_tlast  : out STD_LOGIC;   )           m_axis_tready : in  STD_LOGIC;       =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);   )           s_axis_tvalid : in  STD_LOGIC;   )           s_axis_tlast  : in  STD_LOGIC;   )           s_axis_tready : out STD_LOGIC;�         r      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �  �      �   #        ����                                                                                                                                                                                                                                                                                                                            #           -           V        ^0�     �   "   #          $    signal spi_mosi_tb  : STD_LOGIC;   $    signal spi_miso_tb  : STD_LOGIC;   $    signal stop_data_tb : STD_LOGIC;   +    signal cs_tb        : std_logic := '1';   F    signal outData_tb   : std_logic_vector (7 downto 0) := "01010101";   F    signal inData_tb    : std_logic_vector (7 downto 0) := "00000000";   8    signal ledsData_tb  : std_logic_vector (3 downto 0);   +    signal spi_clk_tb   : STD_LOGIC := '0';   +    signal sys_clk_tb   : STD_LOGIC := '0';   $    signal rst_tb       : STD_LOGIC;   "    signal ii           : integer;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �         g      D           signal m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �         g      0           signal m_axis_tvalid : out STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �         g      0           signal m_axis_tlast  : out STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �         g      0           signal m_axis_tready : in  STD_LOGIC;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �          g      D           signal s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �      !   g      0           signal s_axis_tvalid : in  STD_LOGIC;5�_�  �  �          �   !       ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �       "   g      0           signal s_axis_tlast  : in  STD_LOGIC;5�_�  �  �          �   "       ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �   !   #   g      0           signal s_axis_tready : out STD_LOGIC;5�_�  �  �          �      %    ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �      #   g   	   G           signal m_axis_tdata_tb  : out STD_LOGIC_VECTOR (7 downto 0);   3           signal m_axis_tvalid_tb : out STD_LOGIC;   3           signal m_axis_tlast_tb  : out STD_LOGIC;   3           signal m_axis_tready_tb : in  STD_LOGIC;       G           signal s_axis_tdata_tb  : in  STD_LOGIC_VECTOR (7 downto 0);   3           signal s_axis_tvalid_tb : in  STD_LOGIC;   3           signal s_axis_tlast_tb  : in  STD_LOGIC;   3           signal s_axis_tready_tb : out STD_LOGIC;5�_�  �  �          �   $       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   #   $          D    signal mosiData_tb  : std_logic_vector (7 downto 0):="00000000";5�_�  �  �          �   &       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   %   '   f      7   sys_clk_tb   <= not sys_clk_tb after 100 ns; --10Mhz5�_�  �  �          �   &       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   %   '   f      6   ys_clk_tb   <= not sys_clk_tb after 100 ns; --10Mhz5�_�  �  �          �   &       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   %   '   f      5   s_clk_tb   <= not sys_clk_tb after 100 ns; --10Mhz5�_�  �  �          �   &       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   %   '   f      4   _clk_tb   <= not sys_clk_tb after 100 ns; --10Mhz5�_�  �  �          �   '       ����                                                                                                                                                                                                                                                                                                                               %       "   (          (    ^0�     �   &   (   f         rst_tb   <= '0';5�_�  �             �   (        ����                                                                                                                                                                                                                                                                                                                            (          *           V       ^0�     �   '   (          (--   cs_tb    <= not cs_tb after 320 ns;                   --'0' after 5 ns;    5�_�  �                +        ����                                                                                                                                                                                                                                                                                                                            +           6           V        ^0�     �   *   +                spi_clk_tb <= '1';         cs_tb      <= '1';         wait for 100 ns;         cs_tb<='0';         wait for 100 ns;   (      spi_clk_loop:for k in 0 to 15 loop            wait for 100 ns;   &         spi_clk_tb <= not spi_clk_tb;         end loop spi_clk_loop;         wait for 100 ns;         cs_tb <= '1';         wait for 1000 ns;5�_�                  )        ����                                                                                                                                                                                                                                                                                                                            )          F          V       ^0�     �   (   )             cs_proc: process is      begin      end process;           spi_proc: process(spi_clk_tb)   .      variable i              :integer   := 0;   .      variable inData_integer :integer   := 0;   0      variable mosiData_integer :integer := 100;             begin   *         if falling_edge(spi_clk_tb)  then               if cs_tb = '0' then                  i:=i+1;   -               spi_mosi_tb <= mosiData_tb(7);                  if(i/=8) then   ?                  mosiData_tb <= mosiData_tb(6 downto 0) & '0';                  else   (                  i                := 0;   9                  mosiData_integer := mosiData_integer+1;   j                  mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));   7                  inData_integer   := inData_integer+1;   f                  inData_tb        <= std_logic_vector (to_unsigned(inData_integer,inData_tb'length));                  end if;               else                   i:=0;   g               mosiData_tb      <= std_logic_vector (to_unsigned(mosiData_integer,mosiData_tb'length));               end if;            end if;         ii<=i;      end process;5�_�                 )        ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^0�     �   (   )           5�_�                 +       ����                                                                                                                                                                                                                                                                                                                            +          6                 ^1     �   *   8   8      <           m_axis_tdata   out STD_LOGIC_VECTOR (7 downto 0),   (           m_axis_tvalid  out STD_LOGIC,   (           m_axis_tlast   out STD_LOGIC,   (           m_axis_tready  in  STD_LOGIC,       <           s_axis_tdata   in  STD_LOGIC_VECTOR (7 downto 0),   (           s_axis_tvalid  in  STD_LOGIC,   (           s_axis_tlast   in  STD_LOGIC,   (           s_axis_tready  out STD_LOGIC,       (           clk            in  STD_LOGIC,   )           rst            in  STD_LOGIC),    �   +   ,   8    �   *   7   8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0),   )           m_axis_tvalid : out STD_LOGIC,   )           m_axis_tlast  : out STD_LOGIC,   )           m_axis_tready : in  STD_LOGIC,       =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0),   )           s_axis_tvalid : in  STD_LOGIC,   )           s_axis_tlast  : in  STD_LOGIC,   )           s_axis_tready : out STD_LOGIC,       )           clk           : in  STD_LOGIC,   *           rst           : in  STD_LOGIC),5�_�                 +       ����                                                                                                                                                                                                                                                                                                                            +          6                 ^1
     �   +   7   8      5           m_axis_tvalid m_axis_tvalid out STD_LOGIC,   5           m_axis_tlast  m_axis_tlast  out STD_LOGIC,   5           m_axis_tready m_axis_tready in  STD_LOGIC,   &                                         I           s_axis_tdata  s_axis_tdata  in  STD_LOGIC_VECTOR (7 downto 0),   5           s_axis_tvalid s_axis_tvalid in  STD_LOGIC,   5           s_axis_tlast  s_axis_tlast  in  STD_LOGIC,   5           s_axis_tready s_axis_tready out STD_LOGIC,   &                                         5           clk           clk           in  STD_LOGIC,   6           rst           rst           in  STD_LOGIC),�   *   ,   8      I           m_axis_tdata  m_axis_tdata  out STD_LOGIC_VECTOR (7 downto 0),5�_�                 +   )    ����                                                                                                                                                                                                                                                                                                                            +   )       6   8       ���    ^1     �   *   ,   8      )           m_axis_tdata  =>m_axis_tdata  �   *   7   8      K           m_axis_tdata  =>m_axis_tdata  out STD_LOGIC_VECTOR (7 downto 0),   7           m_axis_tvalid =>m_axis_tvalid out STD_LOGIC,   7           m_axis_tlast  =>m_axis_tlast  out STD_LOGIC,   7           m_axis_tready =>m_axis_tready in  STD_LOGIC,   (                         =>                K           s_axis_tdata  =>s_axis_tdata  in  STD_LOGIC_VECTOR (7 downto 0),   7           s_axis_tvalid =>s_axis_tvalid in  STD_LOGIC,   7           s_axis_tlast  =>s_axis_tlast  in  STD_LOGIC,   7           s_axis_tready =>s_axis_tready out STD_LOGIC,   (                         =>                7           clk           =>clk           in  STD_LOGIC,   8           rst           =>rst           in  STD_LOGIC),5�_�                 6   )    ����                                                                                                                                                                                                                                                                                                                            +   )       6   8       ���    ^1"     �   5   7   8      *           rst           =>rst           ,5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            +   )       6   8       ���    ^1&     �   3   4          (                         =>             5�_�    	             /       ����                                                                                                                                                                                                                                                                                                                            +   )       5   8       ���    ^1(     �   .   /          (                         =>             5�_�    
          	   +   '    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^10     �   *   ,   6      *           m_axis_tdata  =>m_axis_tdata  ,5�_�  	            
   ,   (    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^14     �   +   -   6      *           m_axis_tvalid =>m_axis_tvalid ,5�_�  
               -   '    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^16     �   ,   .   6      *           m_axis_tlast  =>m_axis_tlast  ,5�_�                 .   (    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^17     �   -   /   6      *           m_axis_tready =>m_axis_tready ,5�_�                 /   '    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^18     �   .   0   6      *           s_axis_tdata  =>s_axis_tdata  ,5�_�                 0   (    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^19     �   /   1   6      *           s_axis_tvalid =>s_axis_tvalid ,5�_�                 1   '    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^1:     �   0   2   6      *           s_axis_tlast  =>s_axis_tlast  ,5�_�                 2   (    ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^1;     �   1   3   6      *           s_axis_tready =>s_axis_tready ,5�_�                 3       ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^1=     �   2   4   6      *           clk           =>clk           ,5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            +   )       4   8       ���    ^1?     �   3   5   6      +           rst           =>rst           ),5�_�                 #        ����                                                                                                                                                                                                                                                                                                                                                  V        ^1N     �   "   %   6    �   #   $   6    5�_�                 #       ����                                                                                                                                                                                                                                                                                                                            #          $                 ^1P     �   #   %   8      *           rst           : in  STD_LOGIC);�   "   $   8      )           clk           : in  STD_LOGIC;5�_�                 #       ����                                                                                                                                                                                                                                                                                                                            #          $                 ^1V     �   #   %   8      1           signal rst           : in  STD_LOGIC);�   "   $   8      0           signal clk           : in  STD_LOGIC;5�_�                 #   %    ����                                                                                                                                                                                                                                                                                                                            #   %       $   (          (    ^1Z     �   "   %   8      3           signal clk_tb           : in  STD_LOGIC;   4           signal rst_tb           : in  STD_LOGIC);5�_�                 $   .    ����                                                                                                                                                                                                                                                                                                                            #   %       $   (          (    ^1]     �   #   %   8      0           signal rst_tb           : STD_LOGIC);5�_�                 &       ����                                                                                                                                                                                                                                                                                                                            #   %       $   (          (    ^1_     �   %   '   8            5�_�                 &       ����                                                                                                                                                                                                                                                                                                                            #   %       $   (          (    ^1`     �   %   '   8           5�_�                 &       ����                                                                                                                                                                                                                                                                                                                            #   %       $   (          (    ^1a   w �   %   &              5�_�                 5   -    ����                                                                                                                                                                                                                                                                                                                                                             ^1�   x �   4   6   7      .           rst           =>rst_tb           ),5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             ^1�     �   &   (   7      3   clk_tb   <= not sys_clk_tb after 100 ns; --10Mhz5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             ^1�     �   &   (   7      2   clk_tb   <= not ys_clk_tb after 100 ns; --10Mhz5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                                             ^1�     �   &   (   7      1   clk_tb   <= not s_clk_tb after 100 ns; --10Mhz5�_�                  '       ����                                                                                                                                                                                                                                                                                                                                                             ^1�   y �   &   (   7      0   clk_tb   <= not _clk_tb after 100 ns; --10Mhz5�_�    #                 	    ����                                                                                                                                                                                                                                                                                                                                                             ^1�     �   
      7          port(  5�_�     $  !      #           ����                                                                                                                                                                                                                                                                                                                                      $          V       ^2   { �   #   %          /           signal rst_tb           : STD_LOGIC;�   "   $          /           signal clk_tb           : STD_LOGIC;�   !   #          /           signal s_axis_tready_tb : STD_LOGIC;�       "          /           signal s_axis_tlast_tb  : STD_LOGIC;�      !          /           signal s_axis_tvalid_tb : STD_LOGIC;�                 C           signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0);�                /           signal m_axis_tready_tb : STD_LOGIC;�                /           signal m_axis_tlast_tb  : STD_LOGIC;�                /           signal m_axis_tvalid_tb : STD_LOGIC;�                C           signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0);5�_�  #  %          $   '       ����                                                                                                                                                                                                                                                                                                                                                             ^3�     �   &   (   7    �   '   (   7    5�_�  $  &          %   '       ����                                                                                                                                                                                                                                                                                                                                                             ^3�   | �   &   (   8         rst_tb   <= '0' after 10 ns;5�_�  %  '          &   #   &    ����                                                                                                                                                                                                                                                                                                                                                             ^4     �   "   $   8      '   signal clk_tb           : STD_LOGIC;5�_�  &  (          '   '       ����                                                                                                                                                                                                                                                                                                                                                             ^4   } �   &   '             clk_tb   <= '0' after 10 ns;5�_�  '  )          (   (       ����                                                                                                                                                                                                                                                                                                                                                             ^47     �   (   -   8         �   (   *   7    5�_�  (  *          )   +       ����                                                                                                                                                                                                                                                                                                                                                             ^4L     �   +   -   <            �   +   -   ;    5�_�  )  +          *   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^4R     �   +   -   <            if(ris5�_�  *  ,          +   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^4S     �   +   .   <            if ris5�_�  +  -          ,      :    ����                                                                                                                                                                                                                                                                                                                                                             ^4l     �          =      ;   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0);5�_�  ,  .          -       &    ����                                                                                                                                                                                                                                                                                                                                                             ^4v     �      !   =      '   signal s_axis_tvalid_tb : STD_LOGIC;5�_�  -  /          .       (    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �      !   =      )   signal s_axis_tvalid_tb : STD_LOGIC:=;5�_�  .  0          /       (    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �      !   =      *   signal s_axis_tvalid_tb : STD_LOGIC:=1;5�_�  /  1          0       *    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �      !   =      +   signal s_axis_tvalid_tb : STD_LOGIC:='1;5�_�  0  2          1   !   &    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �       "   =      '   signal s_axis_tlast_tb  : STD_LOGIC;5�_�  1  3          2   "   &    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   !   #   =      '   signal s_axis_tready_tb : STD_LOGIC;5�_�  2  4          3   #   &    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   "   $   =      -   signal clk_tb           : STD_LOGIC :='0';5�_�  3  5          4   $   &    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   #   %   =      '   signal rst_tb           : STD_LOGIC;5�_�  4  6          5   (       ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   '   )   =         rst_tb   <= '0' after 10 ns;5�_�  5  7          6   (       ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   '   )   =         rst_tb   <= '0' after 20 ns;5�_�  6  8          7   (       ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �   '   )   =          rst_tb   <= '0' after 200 ns;5�_�  7  9          8      &    ����                                                                                                                                                                                                                                                                                                                                                             ^4�     �         =      '   signal m_axis_tready_tb : STD_LOGIC;5�_�  8  <          9      &    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^4�     �         =      '   signal m_axis_tready_tb : STD_LOGIC;5�_�  9  =  :      <      &    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^4�   ~ �         =      '   signal m_axis_tlast_tb  : STD_LOGIC;   '   signal m_axis_tready_tb : STD_LOGIC;�         =      '   signal m_axis_tvalid_tb : STD_LOGIC;5�_�  <  >          =   ,       ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5   � �   ,   .   >      	         �   ,   .   =    5�_�  =  ?          >      <    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5A     �          >      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):='01010101';5�_�  >  @          ?      <    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5O     �          >      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):='01010101';5�_�  ?  A          @      E    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5Q   � �          >      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01010101';5�_�  @  C          A   *       ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5X     �   )   +   >         test_proc:process(clk) is5�_�  A  D  B      C   ,       ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5_   � �   +   -   >            if rising_edge(clk) then5�_�  C  E          D      )    ����                                                                                                                                                                :                                                                                                                                                             &          &          &    ^:;   � �         >      ,   signal m_axis_tready_tb : STD_LOGIC:='0';5�_�  D  F          E   (       ����                                                                                                                                                                :                                                                                                                                                             &          &          &    ^:�   � �   '   )   >          rst_tb   <= '0' after 180 ns;5�_�  E  G          F   $   )    ����                                                                                                                                                                :                                                                                                                                                             &          &          &    ^:�   � �   #   %   >      ,   signal rst_tb           : STD_LOGIC:='1';5�_�  F  H          G      :    ����                                                                                                                                                                :                                                                                                                                                             &          &          &    ^;   � �         >      ;   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0);5�_�  G  I          H      ?    ����                                                                                                                                                                :                                                                                                                                                             
                 v       ^;}     �          >      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01010101";5�_�  H  J          I      C    ����                                                                                                                                                                :                                                                                                                                                             
                 v       ^;~   � �          >      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110101";5�_�  I  K          J   *       ����                                                                                                                                                                :                                                                                                                                                             
                 v       ^I�     �   )   +   >         test_proc:process(clk_tb) is5�_�  J  L          K   ,       ����                                                                                                                                                                :                                                                                                                                                             
                 v       ^I�     �   +   -   >      !      if rising_edge(clk_tb) then5�_�  K  M          L   ,   !    ����                                                                                                                                                                :                                                                                                                                                             
                 v       ^I�     �   ,   .   >    5�_�  L  N          M      
    ����                                                                                                                                                                ;                                                                                                                                                             
                 v       ^I�     �          ?      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";5�_�  M  O          N   -        ����                                                                                                                                                                ;                                                                                                                                                             
                 v       ^I�     �   ,   .   ?       �   -   .   ?    5�_�  N  P          O   -        ����                                                                                                                                                                ;                                                                                                                                                          -          -          V   
    ^I�     �   ,   .   >    �   -   .   >    �   ,   -          clk_tb5�_�  O  Q          P   -        ����                                                                                                                                                                ;                                                                                                                                                          -           -          V   
    ^I�     �   ,   .          s_axis_tdata_tb5�_�  P  R          Q   -       ����                                                                                                                                                                ;                                                                                                                                                          -           -          V   
    ^I�   � �   ,   .   ?               s_axis_tdata_tb5�_�  Q  T          R   *   "    ����                                                                                                                                                                ;                                                                                                                                                          -           -          V   
    ^I�     �   )   +   ?      &   test_proc:process(s_axis_tready) is5�_�  R  U  S      T   ,   "    ����                                                                                                                                                                ;                                                                                                                                                          -           -          V   
    ^I�   � �   +   -   ?      (      if rising_edge(s_axis_tready) then5�_�  T  V          U   2        ����                                                                                                                                                                ;                                                                                                                                                                                           ^�     �   1   3   ?      stretcher_inst:stretcher5�_�  U  W          V   2       ����                                                                                                                                                                ;                                                                                                                                                                                           ^�*     �   1   3   ?      split_8to1_inst:stretcher5�_�  V  X          W   
       ����                                                                                                                                                                ;                                                                                                                                                                                           ^�7     �   	      ?         component stretcher is5�_�  W  Y          X          ����                                                                                                                                                                ;                                                                                                                                                                                           ^�:   � �         ?         end component stretcher;5�_�  X  Z          Y   
        ����                                                                                                                                                                ;                                                                                                                                                                                           ^�j   � �   1   3          split_8to1_inst:split_8to1�                   end component split_8to1;�   	                component split_8to1 is5�_�  Y              Z           ����                                                                                                                                                                :                                                                                                                                                                                           ^Y     �              �          >       5�_�  R          T  S   ,   #    ����                                                                                                                                                                ;                                                                                                                                                          -           -          V   
    ^I�     �   +   -   ?      +      if rising_edge(s_axis_tready)_tb then5�_�  A          C  B   ,       ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^5\     �   +   -   >      !      if rising_edge(clk)_tb then5�_�  9  ;      <  :      &    ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^4�     �         =      (   signal m_axis_tvalid_tb : STD_LOGIC:;5�_�  :              ;          ����                                                                                                                                                                                                                                                                                                                               &          &          &    ^4�     �         =         end component stretcher;=5�_�     "      #  !          ����                                                                                                                                                                                                                                                                                                                                                             ^1�     �         7         end componentstretcher;5�_�  !              "          ����                                                                                                                                                                                                                                                                                                                                                             ^1�   z �         7         end component;5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                            #           #           V        ^0�     �         g      3           signal m_axis_tvali_tbd : out STD_LOGIC;5�_�  �          �  �   #        ����                                                                                                                                                                                                                                                                                                                            #          #          V       ^0�     �   "   ,        5�_�  �          �  �   ;       ����                                                                                                                                                                                                                                                                                                                                                             ^/�     �   :   <   c      )   stretcherspi_proc: process(spi_clk_tb)5�_�  �  �      �  �   %       ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      -   pi_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �  �          �   %       ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      ,   i_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �              �   %       ����                                                                                                                                                                                                                                                                                                                                                        ^J�     �   $   &   c      ,   c_clk_tb   <= not spi_clk_tb after 20 ns;5�_�  �          �  �   T       ����                                                                                                                                                                                                                                                                                                                            *   
       +   
       V   
    ^B9     �   S   U   _       5�_�  T          V  U   -   	    ����                                                                                                                                                                                                                                                                                                                            /          9          V       ^�Q     �   ,   .        5�_�                 F        ����                                                                                                                                                                                                                                                                                                                            @          @   %       v   %    ^�m   I �   E   G          fnd arq;5�_�  
                      ����                                                                                                                                                                                                                                                                                                                            )          )          V       ]��B     �         F      7    ignal mosiData_tb  : std_logic_vector (7 downto 0);5�_�                +   !    ����                                                                                                                                                                                                                                                                                                                            0          1          V       ]���     �   *   ,   D      ,         spi_mosi_tb <= mosiData_integer(7);5�_�                   -   &    ����                                                                                                                                                                                                                                                                                                                            0          1          V       ]���   ? �   ,   .   D      @            mosiData_tb   <= mosiData_integer(6 downto 0) & '0';5�_�   �           �   �   *        ����                                                                                                                                                                                                                                                                                                                            *           0           V        ]��3     �   )   +          &         spi_mosi_tb <= outData_tb(7);�   +   -          9            outData_tb   <= outData_tb(6 downto 0) & '0';�   .   0          1            outData_integer := outData_integer+1;�   /   1          a            outData_tb      <= std_logic_vector (to_unsigned(outData_integer,outData_tb'length));5�_�   �       �   �   �   8        ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�,s     �   7   ?   A      (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   8        ����                                                                                                                                                                                                                                                                                                                            8          >          V       ]�,p     �   7   ?   A      (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   ,eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   0   H    ����                                                                                                                                                                                                                                                                                                                            0   H       0   \       v   \    ]�     �   /   1   @      O            inData_tb   <= std_logic_vector (to_unsigned(inData_integer,) + 1);5�_�   �           �   �   %        ����                                                                                                                                                                                                                                                                                                                            %           &           V        ]�Z     �   $   '   A      )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   %       ����                                                                                                                                                                                                                                                                                                                            &          %          V       ]�S     �   $   '   A      eeeeeeeeeeeeeeeeeeeeeeeeeee   (eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                            .   	       0   	       V   	    ]�#     �         @      K    signal inData_tb_shift   : std_logic_vector (7 downto 0) := "00000000";5�_�   �           �   �   ,        ����                                                                                                                                                                                                                                                                                                                            "   	       "   	       V   	    ]��     �   ,   -   <    �   ,   -   <         loop_proc: process      variable i: integer := 0;      begin         for i in 0 to 10 loop            wait for 320 ns;   A         inData_tb <= std_logic_vector (unsigned(inData_tb) + 1);         end loop;      end process;5�_�   �           �   �   -       ����                                                                                                                                                                                                                                                                                                                            1          1          V       ]��     �   ,   .   >      "      if(rising_edge(clk)_tb) then5�_�   �           �   �   .   1    ����                                                                                                                                                                                                                                                                                                                            "          )          V       ]��     �   .   /   C      	         �   .   0   D               endifh5�_�   7   9       :   8           ����                                                                                                                                                                                                                                                                                                                                                V       ]��B     �              5�_�   8               9           ����                                                                                                                                                                                                                                                                                                                                                V       ]��D    �             �               )    signal spi_mosi_tb : in    STD_LOGIC;   )    signal spi_miso_tb : out   STD_LOGIC;   )    signal cs_tb       : in    std_logic;   =    signal outData_tb  : out   std_logic_vector (7 downto 0);   =    signal inData_tb   : in    std_logic_vector (7 downto 0);   =    signal ledsData_tb : out   std_logic_vector (3 downto 0);   )    signal clk_tb      : in    STD_LOGIC;5�_�   '           )   (   ?   #    ����                                                                                                                                                                                                                                                                                                                            :   #       ?   #          #    ]���     �   >   @   B      ,           ledsData     => ledsDatakkkkkkk ,5�_�                    :        ����                                                                                                                                                                                                                                                                                                                            :   )       @   %       V   )    ]��v     �   9   A   C      *eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   :eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   :eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   :eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   %eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�                    :        ����                                                                                                                                                                                                                                                                                                                            :           A   	       V        ]��_     �   9   ;        �   :   ;        �   9   :   :      &    port ( spi_mosi : in    STD_LOGIC;   &           spi_miso : out   STD_LOGIC;   &           cs       : in    std_logic;   :           outData  : out   std_logic_vector (7 downto 0);   :           inData   : in    std_logic_vector (7 downto 0);   :           ledsData : out   std_logic_vector (3 downto 0);   %           clk      : in    STD_LOGIC   
        );5��