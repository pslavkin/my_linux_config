Vim�UnDo� �ӕRs����5���'7Kt���ʱ����E  ?                '      '  '  '    ^$G�   � _�                     1        ����                                                                                                                                                                                                                                                                                                                                                             ^�W     �   0   U   ?    �   1   2   ?    5�_�                    1       ����                                                                                                                                                                                                                                                                                                                                                             ^�X     �   0   2   c         shift_reg:process (clk) is5�_�                    0   
    ����                                                                                                                                                                                                                                                                                                                                                             ^�]     �   0   2   c    5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             ^�`     �   1   3   d         axi_proc:process (clk) is5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                                             ^�     �         d    �   	   
   d    5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �      
   f      5   type shiftState is (waitingSvalid, waitingMready);5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   	      f      ,   signal state:shiftState := waitingSvalid;5�_�      	              1        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   0   1           5�_�      
           	   0       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   /   1                   end if;5�_�   	              
   9       ����                                                                                                                                                                                                                                                                                                                            9          :                 ^��     �   9   ;   e      !            m_axis_tvalid <= '0';�   8   :   e      !            s_axis_tready <= '1';5�_�   
                 ;       ����                                                                                                                                                                                                                                                                                                                            9          :                 ^��     �   :   <   e      -            m_axis_tdata  <= (others => '0');5�_�                    ?   "    ����                                                                                                                                                                                                                                                                                                                            ?   "       @   "          "    ^��     �   ?   A   e      ,                     s_axis_tready   <= '0';�   >   @   e      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo5�_�                    B   !    ����                                                                                                                                                                                                                                                                                                                            B   !       C   !          !    ^��     �   B   D   e      V                     m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato�   A   C   e      T                     m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    D   "    ����                                                                                                                                                                                                                                                                                                                            B   !       C   !          !    ^��     �   C   E   e      q                     m_axis_tvalid   <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�                    E   %    ����                                                                                                                                                                                                                                                                                                                            B   !       C   !          !    ^��     �   D   F   e                           state           <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato5�_�                    B   7    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   B   D   e      Y                     m_axis_tdata_tb(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato�   A   C   e      W                     m_axis_tdata_tb(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    H   "    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   G   I   e      q                  if m_axis_tready = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�                   K   $    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   J   L   e      W                        m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    L   $    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   K   M   e      Y                        m_axis_tdata(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�                    K   :    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   J   L   e      Z                        m_axis_tdata_tb(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                    L   :    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   K   M   e      \                        m_axis_tdata_tb(1) <= s_axis_tdata(bitCounter+1);    --pongo el dato5�_�                    N   %    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   M   O   e      �                        m_axis_tvalid <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�                    O   %    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   N   P   e      -                        s_axis_tready <= '1';5�_�                    V       ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��    �   U   W   e         end process shift_reg;5�_�                   9       ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^M     �   8   :   e    �   9   :   e    5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            C   7       D   7          7    ^P     �   9   ;   f      $            s_axis_tready_tb <= '1';5�_�                    :   !    ����                                                                                                                                                                                                                                                                                                                            C   7       D   7          7    ^R     �   9   ;   f      !            s_axis_tvalid <= '1';5�_�                    9        ����                                                                                                                                                                                                                                                                                                                            9   #       <   0       V   P    ^`     �   c   e   f      .           rst           =>rst_tb           );�   b   d   f      -           clk           =>clk_tb           ,�   a   c   f      -           s_axis_tready =>s_axis_tready_tb ,�   `   b   f      -           s_axis_tlast  =>s_axis_tlast_tb  ,�   _   a   f      -           s_axis_tvalid =>s_axis_tvalid_tb ,�   ^   `   f      -           s_axis_tdata  =>s_axis_tdata_tb  ,�   ]   _   f      -           m_axis_tready =>m_axis_tready_tb ,�   \   ^   f      -           m_axis_tlast  =>m_axis_tlast_tb  ,�   [   ]   f      -           m_axis_tvalid =>m_axis_tvalid_tb ,�   Z   \   f      -           m_axis_tdata  =>m_axis_tdata_tb  ,�   Y   [   f          port map(  �   V   X   f         end process axi_master_proc;�   U   W   f            end if;�   T   V   f               end if;�   S   U   f                  end case;�   R   T   f                        end if;�   Q   S   f                           end if;�   P   R   f      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   O   Q   f      0                        s_axis_tready_tb <= '1';�   N   P   f      �                        m_axis_tvalid_tb <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   M   O   f                           else�   L   N   f      _                        m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   K   M   f      ]                        m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   J   L   f      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   I   K   f      Q                     bitCounter := bitCounter+2;                     --incremento�   H   J   f      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   G   I   f      $               when waitingMready =>�   F   H   f                        end if;�   E   G   f      �                     state              <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   D   F   f      t                     m_axis_tvalid_tb   <= '1';                         --como puedo mandar, le avoso que tengo dato�   C   E   f      \                     m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   B   D   f      Z                     m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   A   C   f      *                     bitCounter      := 0;�   @   B   f      /                     s_axis_tready_tb   <= '0';�   ?   A   f      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   >   @   f      $               when waitingSvalid =>�   =   ?   f                  case state is�   <   >   f               else�   ;   =   f      0            m_axis_tdata_tb  <= (others => '0');�   :   <   f      $            m_axis_tvalid_tb <= '0';�   9   ;   f      T            s_axis_tvalid    <= '1'; --que haga de cuentqa que siempre tiene un dato�   8   :   f      $            s_axis_tready_tb <= '1';�   7   9   f      +            state         <= waitingSvalid;�   6   8   f               if rst = '0' then�   5   7   f            if rising_edge(clk) then�   4   6   f         begin�   3   5   f      0      variable bitCounter :integer range 0 to 8;�   2   4   f      #   axi_master_proc:process (clk) is�   0   2   f         end process test_proc;�   /   1   f            end if;�   .   0   f      '         s_axis_tdata_tb <= "10010101";�   -   /   f      +      if rising_edge(s_axis_tready_tb) then�   ,   .   f         begin�   +   -   f      )   test_proc:process(s_axis_tready_tb) is�   )   +   f          rst_tb   <= '1' after 180 ns;�   (   *   f      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   %   '   f      ,   signal rst_tb           : STD_LOGIC:='0';�   $   &   f      ,   signal clk_tb           : STD_LOGIC:='0';�   #   %   f      ,   signal s_axis_tready_tb : STD_LOGIC:='0';�   "   $   f      ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';�   !   #   f      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';�       "   f      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";�          f      ,   signal m_axis_tready_tb : STD_LOGIC:='1';�         f      ,   signal m_axis_tlast_tb  : STD_LOGIC:='0';�         f      ,   signal m_axis_tvalid_tb : STD_LOGIC:='0';�         f      J   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         f         end component split_1to8;�         f      *           rst           : in  STD_LOGIC);�         f      )           clk           : in  STD_LOGIC;�         f      )           s_axis_tready : out STD_LOGIC;�         f      )           s_axis_tlast  : in  STD_LOGIC;�         f      )           s_axis_tvalid : in  STD_LOGIC;�         f      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         f      )           m_axis_tready : in  STD_LOGIC;�         f      )           m_axis_tlast  : out STD_LOGIC;�         f      )           m_axis_tvalid : out STD_LOGIC;�         f      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         f      	    port(�         f         component split_1to8 is�   	      f      +   signal state:axiStates := waitingSvalid;�      
   f      4   type axiStates is (waitingSvalid, waitingMready);�   8   :          $            s_axis_tready_tb <= '1';�   ;   =          0            m_axis_tdata_tb  <= (others => '0');�   :   <          $            m_axis_tvalid_tb <= '0';�   9   ;          Q            s_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�                     A        ����                                                                                                                                                                                                                                                                                                                            A   &       F   &       V   &    ^v     �   c   e   f      .           rst           =>rst_tb           );�   b   d   f      -           clk           =>clk_tb           ,�   a   c   f      -           s_axis_tready =>s_axis_tready_tb ,�   `   b   f      -           s_axis_tlast  =>s_axis_tlast_tb  ,�   _   a   f      -           s_axis_tvalid =>s_axis_tvalid_tb ,�   ^   `   f      -           s_axis_tdata  =>s_axis_tdata_tb  ,�   ]   _   f      -           m_axis_tready =>m_axis_tready_tb ,�   \   ^   f      -           m_axis_tlast  =>m_axis_tlast_tb  ,�   [   ]   f      -           m_axis_tvalid =>m_axis_tvalid_tb ,�   Z   \   f      -           m_axis_tdata  =>m_axis_tdata_tb  ,�   Y   [   f          port map(  �   V   X   f         end process axi_master_proc;�   U   W   f            end if;�   T   V   f               end if;�   S   U   f                  end case;�   R   T   f                        end if;�   Q   S   f                           end if;�   P   R   f      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   O   Q   f      0                        s_axis_tready_tb <= '1';�   N   P   f      �                        m_axis_tvalid_tb <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   M   O   f                           else�   L   N   f      _                        m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   K   M   f      ]                        m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   J   L   f      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   I   K   f      Q                     bitCounter := bitCounter+2;                     --incremento�   H   J   f      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   G   I   f      $               when waitingMready =>�   F   H   f                        end if;�   E   G   f      �                     state              <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   D   F   f      t                     m_axis_tvalid_tb   <= '1';                         --como puedo mandar, le avoso que tengo dato�   C   E   f      \                     m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   B   D   f      Z                     m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   A   C   f      -                     bitCounter         := 0;�   @   B   f      /                     s_axis_tready_tb   <= '0';�   ?   A   f      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   >   @   f      $               when waitingSvalid =>�   =   ?   f                  case state is�   <   >   f               else�   ;   =   f      0            m_axis_tdata_tb  <= (others => '0');�   :   <   f      $            m_axis_tvalid_tb <= '0';�   9   ;   f      T            s_axis_tvalid    <= '1'; --que haga de cuentqa que siempre tiene un dato�   8   :   f      $            s_axis_tready_tb <= '1';�   7   9   f      +            state         <= waitingSvalid;�   6   8   f               if rst = '0' then�   5   7   f            if rising_edge(clk) then�   4   6   f         begin�   3   5   f      0      variable bitCounter :integer range 0 to 8;�   2   4   f      #   axi_master_proc:process (clk) is�   0   2   f         end process test_proc;�   /   1   f            end if;�   .   0   f      '         s_axis_tdata_tb <= "10010101";�   -   /   f      +      if rising_edge(s_axis_tready_tb) then�   ,   .   f         begin�   +   -   f      )   test_proc:process(s_axis_tready_tb) is�   )   +   f          rst_tb   <= '1' after 180 ns;�   (   *   f      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   %   '   f      ,   signal rst_tb           : STD_LOGIC:='0';�   $   &   f      ,   signal clk_tb           : STD_LOGIC:='0';�   #   %   f      ,   signal s_axis_tready_tb : STD_LOGIC:='0';�   "   $   f      ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';�   !   #   f      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';�       "   f      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";�          f      ,   signal m_axis_tready_tb : STD_LOGIC:='1';�         f      ,   signal m_axis_tlast_tb  : STD_LOGIC:='0';�         f      ,   signal m_axis_tvalid_tb : STD_LOGIC:='0';�         f      J   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         f         end component split_1to8;�         f      *           rst           : in  STD_LOGIC);�         f      )           clk           : in  STD_LOGIC;�         f      )           s_axis_tready : out STD_LOGIC;�         f      )           s_axis_tlast  : in  STD_LOGIC;�         f      )           s_axis_tvalid : in  STD_LOGIC;�         f      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         f      )           m_axis_tready : in  STD_LOGIC;�         f      )           m_axis_tlast  : out STD_LOGIC;�         f      )           m_axis_tvalid : out STD_LOGIC;�         f      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         f      	    port(�         f         component split_1to8 is�   	      f      +   signal state:axiStates := waitingSvalid;�      
   f      4   type axiStates is (waitingSvalid, waitingMready);�   @   B          /                     s_axis_tready_tb   <= '0';�   E   G          �                     state              <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   D   F          t                     m_axis_tvalid_tb   <= '1';                         --como puedo mandar, le avoso que tengo dato�   C   E          \                     m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   B   D          Z                     m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   A   C          *                     bitCounter      := 0;5�_�      !               C   $    ����                                                                                                                                                                                                                                                                                                                            A   &       F   &       V   &    ^{     �   B   D   f      Z                     m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�       "           !   C   $    ����                                                                                                                                                                                                                                                                                                                            A   &       F   &       V   &    ^{     �   B   D   f      Y                     m_axis_tdata_tb0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   !   #           "   C   $    ����                                                                                                                                                                                                                                                                                                                            A   &       F   &       V   &    ^|     �   B   D   f      X                     m_axis_tdata_tb) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   "   $           #   C   (    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^~     �   B   D   f      W                     m_axis_tdata_tb <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   #   %           $   C   (    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   B   D   f      <                     m_axis_tdata_tb <= ;    --pongo el dato5�_�   $   &           %   C   3    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   B   D   f      F                     m_axis_tdata_tb <= "10101100";    --pongo el dato5�_�   %   '           &   D       ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   C   D          \                     m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato5�_�   &   (           '   C   (    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   B   D   e      3                     m_axis_tdata_tb <= "10101100";5�_�   '   )           (   C   F    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   B   D   e      Q                     m_axis_tdata_tb <= STD_LOGIC_VECTOR(signed(data))"10101100";5�_�   (   *           )   4   /    ����                                                                                                                                                                                                                                                                                                                            C   (       C   B       v   B    ^�     �   3   5   e    �   4   5   e    5�_�   )   +           *   5       ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      0      variable bitCounter :integer range 0 to 8;5�_�   *   ,           +   5   #    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      *      variable data :integer range 0 to 8;5�_�   +   -           ,   5   '    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      .      variable data :integer range -1280 to 8;5�_�   ,   .           -   5   +    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      -      variable data :integer range -128 to 8;5�_�   -   /           .   5   -    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      /      variable data :integer range -128 to 128;5�_�   .   0           /   5   -    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      /      variable data :integer range -128 to 128;5�_�   /   1           0   5   .    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   4   6   f      /      variable data :integer range -128 to 127;5�_�   0   2           1   =   /    ����                                                                                                                                                                                                                                                                                                                            D   (       D   B       v   B    ^�     �   <   >   f    �   =   >   f    5�_�   1   3           2   >       ����                                                                                                                                                                                                                                                                                                                            E   (       E   B       v   B    ^�     �   =   ?   g      0            m_axis_tdata_tb  <= (others => '0');5�_�   2   4           3   >       ����                                                                                                                                                                                                                                                                                                                            E   (       E   B       v   B    ^�     �   =   ?   g      %            data  <= (others => '0');5�_�   3   5           4   >       ����                                                                                                                                                                                                                                                                                                                            E   (       E   B       v   B    ^�     �   =   ?   g      %            data  := (others => '0');5�_�   4   6           5   >       ����                                                                                                                                                                                                                                                                                                                            E   (       E   B       v   B    ^�     �   =   ?   g                  data  := ;5�_�   5   7           6   E       ����                                                                                                                                                                                                                                                                                                                            E   (       E   B       v   B    ^�     �   E   G   h                           �   E   G   g    5�_�   6   8           7   C        ����                                                                                                                                                                                                                                                                                                                            C   %       H   %       V   %    ^�     �   e   g   h      .           rst           =>rst_tb           );�   d   f   h      -           clk           =>clk_tb           ,�   c   e   h      -           s_axis_tready =>s_axis_tready_tb ,�   b   d   h      -           s_axis_tlast  =>s_axis_tlast_tb  ,�   a   c   h      -           s_axis_tvalid =>s_axis_tvalid_tb ,�   `   b   h      -           s_axis_tdata  =>s_axis_tdata_tb  ,�   _   a   h      -           m_axis_tready =>m_axis_tready_tb ,�   ^   `   h      -           m_axis_tlast  =>m_axis_tlast_tb  ,�   ]   _   h      -           m_axis_tvalid =>m_axis_tvalid_tb ,�   \   ^   h      -           m_axis_tdata  =>m_axis_tdata_tb  ,�   [   ]   h          port map(  �   X   Z   h         end process axi_master_proc;�   W   Y   h            end if;�   V   X   h               end if;�   U   W   h                  end case;�   T   V   h                        end if;�   S   U   h                           end if;�   R   T   h      �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   Q   S   h      0                        s_axis_tready_tb <= '1';�   P   R   h      �                        m_axis_tvalid_tb <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   O   Q   h                           else�   N   P   h      _                        m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato�   M   O   h      ]                        m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato�   L   N   h      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   �   K   M   h      Q                     bitCounter := bitCounter+2;                     --incremento�   J   L   h      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   I   K   h      $               when waitingMready =>�   H   J   h                        end if;�   G   I   h      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   F   H   h      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   E   G   h      2                     data             := data + 1;�   D   F   h      H                     m_axis_tdata_tb  <= STD_LOGIC_VECTOR(signed(data));�   C   E   h      +                     bitCounter       := 0;�   B   D   h      -                     s_axis_tready_tb <= '0';�   A   C   h      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   @   B   h      $               when waitingSvalid =>�   ?   A   h                  case state is�   >   @   h               else�   =   ?   h                  data  := 0;�   <   >   h      0            m_axis_tdata_tb  <= (others => '0');�   ;   =   h      $            m_axis_tvalid_tb <= '0';�   :   <   h      T            s_axis_tvalid    <= '1'; --que haga de cuentqa que siempre tiene un dato�   9   ;   h      $            s_axis_tready_tb <= '1';�   8   :   h      +            state         <= waitingSvalid;�   7   9   h               if rst = '0' then�   6   8   h            if rising_edge(clk) then�   5   7   h         begin�   4   6   h      2      variable data :integer range -128 to 127:=0;�   3   5   h      0      variable bitCounter :integer range 0 to 8;�   2   4   h      #   axi_master_proc:process (clk) is�   0   2   h         end process test_proc;�   /   1   h            end if;�   .   0   h      '         s_axis_tdata_tb <= "10010101";�   -   /   h      +      if rising_edge(s_axis_tready_tb) then�   ,   .   h         begin�   +   -   h      )   test_proc:process(s_axis_tready_tb) is�   )   +   h          rst_tb   <= '1' after 180 ns;�   (   *   h      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   %   '   h      ,   signal rst_tb           : STD_LOGIC:='0';�   $   &   h      ,   signal clk_tb           : STD_LOGIC:='0';�   #   %   h      ,   signal s_axis_tready_tb : STD_LOGIC:='0';�   "   $   h      ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';�   !   #   h      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';�       "   h      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";�          h      ,   signal m_axis_tready_tb : STD_LOGIC:='1';�         h      ,   signal m_axis_tlast_tb  : STD_LOGIC:='0';�         h      ,   signal m_axis_tvalid_tb : STD_LOGIC:='0';�         h      J   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         h         end component split_1to8;�         h      *           rst           : in  STD_LOGIC);�         h      )           clk           : in  STD_LOGIC;�         h      )           s_axis_tready : out STD_LOGIC;�         h      )           s_axis_tlast  : in  STD_LOGIC;�         h      )           s_axis_tvalid : in  STD_LOGIC;�         h      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         h      )           m_axis_tready : in  STD_LOGIC;�         h      )           m_axis_tlast  : out STD_LOGIC;�         h      )           m_axis_tvalid : out STD_LOGIC;�         h      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         h      	    port(�         h         component split_1to8 is�   	      h      +   signal state:axiStates := waitingSvalid;�      
   h      4   type axiStates is (waitingSvalid, waitingMready);�   B   D          /                     s_axis_tready_tb   <= '0';�   G   I          �                     state              <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   D   F          G                     m_axis_tdata_tb <= STD_LOGIC_VECTOR(signed(data));�   C   E          -                     bitCounter         := 0;�   F   H          t                     m_axis_tvalid_tb   <= '1';                         --como puedo mandar, le avoso que tengo dato�   E   G          &                     data := data + 1;5�_�   7   9           8   E   )    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^      �   D   F   h      H                     m_axis_tdata_tb  <= STD_LOGIC_VECTOR(signed(data));5�_�   8   :           9   L   .    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^	     �   K   M   h      Q                     bitCounter := bitCounter+2;                     --incremento5�_�   9   ;           :   M   %    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^     �   L   N   h      f                     if bitCounter < 8 then                             --perfecto, porque bit voy?   5�_�   :   <           ;   N   '    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^     �   M   O   h      ]                        m_axis_tdata_tb(0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   ;   =           <   N   '    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^     �   M   O   h      \                        m_axis_tdata_tb0) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   <   >           =   N   '    ����                                                                                                                                                                                                                                                                                                                            E   )       E   8       v   8    ^     �   M   O   h      [                        m_axis_tdata_tb) <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   =   ?           >   N        ����                                                                                                                                                                                                                                                                                                                            N   -       N   -       V   -    ^     �   M   O   g    �   N   O   g    �   M   N          Z                        m_axis_tdata_tb <= s_axis_tdata_tb(bitCounter);    --pongo el dato5�_�   >   @           ?   O       ����                                                                                                                                                                                                                                                                                                                            N           N   G       V   -    ^     �   N   O          _                        m_axis_tdata_tb(1) <= s_axis_tdata_tb(bitCounter+1);    --pongo el dato5�_�   ?   A           @   N       ����                                                                                                                                                                                                                                                                                                                            N           N   G       V   -    ^     �   M   O          H                     m_axis_tdata_tb  <= std_logic_vector(signed(data));5�_�   @   B           A   P        ����                                                                                                                                                                                                                                                                                                                            P          R          V       ^     �   d   f   g      .           rst           =>rst_tb           );�   c   e   g      -           clk           =>clk_tb           ,�   b   d   g      -           s_axis_tready =>s_axis_tready_tb ,�   a   c   g      -           s_axis_tlast  =>s_axis_tlast_tb  ,�   `   b   g      -           s_axis_tvalid =>s_axis_tvalid_tb ,�   _   a   g      -           s_axis_tdata  =>s_axis_tdata_tb  ,�   ^   `   g      -           m_axis_tready =>m_axis_tready_tb ,�   ]   _   g      -           m_axis_tlast  =>m_axis_tlast_tb  ,�   \   ^   g      -           m_axis_tvalid =>m_axis_tvalid_tb ,�   [   ]   g      -           m_axis_tdata  =>m_axis_tdata_tb  ,�   Z   \   g          port map(  �   W   Y   g         end process axi_master_proc;�   V   X   g            end if;�   U   W   g               end if;�   T   V   g                  end case;�   S   U   g                        end if;�   R   T   g                           end if;�   Q   S   g      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   P   R   g      0                        s_axis_tready_tb <= '1';�   O   Q   g      �                        m_axis_tvalid_tb <= '0';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   N   P   g                           else�   M   O   g      K                        m_axis_tdata_tb  <= std_logic_vector(signed(data));�   L   N   g      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   K   M   g      Q                     bitCounter := bitCounter+1;                     --incremento�   J   L   g      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   I   K   g      $               when waitingMready =>�   H   J   g                        end if;�   G   I   g      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   F   H   g      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   E   G   g      2                     data             := data + 1;�   D   F   g      H                     m_axis_tdata_tb  <= std_logic_vector(signed(data));�   C   E   g      +                     bitCounter       := 0;�   B   D   g      -                     s_axis_tready_tb <= '0';�   A   C   g      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   @   B   g      $               when waitingSvalid =>�   ?   A   g                  case state is�   >   @   g               else�   =   ?   g                  data  := 0;�   <   >   g      0            m_axis_tdata_tb  <= (others => '0');�   ;   =   g      $            m_axis_tvalid_tb <= '0';�   :   <   g      T            s_axis_tvalid    <= '1'; --que haga de cuentqa que siempre tiene un dato�   9   ;   g      $            s_axis_tready_tb <= '1';�   8   :   g      +            state         <= waitingSvalid;�   7   9   g               if rst = '0' then�   6   8   g            if rising_edge(clk) then�   5   7   g         begin�   4   6   g      2      variable data :integer range -128 to 127:=0;�   3   5   g      0      variable bitCounter :integer range 0 to 8;�   2   4   g      #   axi_master_proc:process (clk) is�   0   2   g         end process test_proc;�   /   1   g            end if;�   .   0   g      '         s_axis_tdata_tb <= "10010101";�   -   /   g      +      if rising_edge(s_axis_tready_tb) then�   ,   .   g         begin�   +   -   g      )   test_proc:process(s_axis_tready_tb) is�   )   +   g          rst_tb   <= '1' after 180 ns;�   (   *   g      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   %   '   g      ,   signal rst_tb           : STD_LOGIC:='0';�   $   &   g      ,   signal clk_tb           : STD_LOGIC:='0';�   #   %   g      ,   signal s_axis_tready_tb : STD_LOGIC:='0';�   "   $   g      ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';�   !   #   g      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';�       "   g      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";�          g      ,   signal m_axis_tready_tb : STD_LOGIC:='1';�         g      ,   signal m_axis_tlast_tb  : STD_LOGIC:='0';�         g      ,   signal m_axis_tvalid_tb : STD_LOGIC:='0';�         g      J   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         g         end component split_1to8;�         g      *           rst           : in  STD_LOGIC);�         g      )           clk           : in  STD_LOGIC;�         g      )           s_axis_tready : out STD_LOGIC;�         g      )           s_axis_tlast  : in  STD_LOGIC;�         g      )           s_axis_tvalid : in  STD_LOGIC;�         g      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         g      )           m_axis_tready : in  STD_LOGIC;�         g      )           m_axis_tlast  : out STD_LOGIC;�         g      )           m_axis_tvalid : out STD_LOGIC;�         g      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         g      	    port(�         g         component split_1to8 is�   	      g      +   signal state:axiStates := waitingSvalid;�      
   g      4   type axiStates is (waitingSvalid, waitingMready);�   O   Q          �                        m_axis_tvalid_tb <= '0' ;                          --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   Q   S          �                        state         <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   P   R          0                        s_axis_tready_tb <= '1';5�_�   A   C           B   P   0    ����                                                                                                                                                                                                                                                                                                                            P          R          V       ^!     �   O   Q   g      �                        m_axis_tvalid_tb <= '0';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�   B   D           C   -        ����                                                                                                                                                                                                                                                                                                                            ,   (       2           V   /    ^1     �   +   -   a      )   test_proc:process(s_axis_tready_tb) is�   ,   -             begin   +      if rising_edge(s_axis_tready_tb) then   '         s_axis_tdata_tb <= "10010101";         end if;      end process test_proc;    5�_�   C   E           D   ,        ����                                                                                                                                                                                                                                                                                                                            ,   (       -           V   /    ^2    �   +   ,           5�_�   D   F           E           ����                                                                                                                                                                                                                                                                                                                                                             ^�    �      	          architecture arq of tp_tb is�                entity tp_tb is5�_�   E   G           F           ����                                                                                                                                                                                                                                                                                                                                                  V        ^�    �         `      use IEEE.NUMERIC_STD.ALL;5�_�   F   I           G   ,       ����                                                                                                                                                                                                                                                                                                                                                             ^L     �   +   -   `      #   axi_master_proc:process (clk) is5�_�   G   J   H       I   0       ����                                                                                                                                                                                                                                                                                                                                                             ^R    �   /   1   `            if rising_edge(clk) then5�_�   I   K           J   1       ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   0   2   `               if rst = '0' then5�_�   J   L           K   4       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   3   5   `      T            s_axis_tvalid    <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   K   M           L   4       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   3   5   `      W            s_axis_tvalid_tb    <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   L   N           M   4       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   3   5   `      V            s_axis_tvalid_tb   <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   M   O           N   4       ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   3   5   `      U            s_axis_tvalid_tb  <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   N   P           O   >   :    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   =   ?   `      H                     m_axis_tdata_tb  <= std_logic_vector(signed(data));5�_�   O   Q           P   >   H    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   =   ?   `      K                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data));5�_�   P   R           Q   >   I    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   =   ?   `      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   Q   S           R   >   T    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   =   ?   `      X                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,data'length8));5�_�   R   T           S   G   J    ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   F   H   `    �   G   H   `    5�_�   S   U           T   H       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   G   H          K                        m_axis_tdata_tb  <= std_logic_vector(signed(data));5�_�   T   W           U   G       ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   F   H          W                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,data'length));5�_�   U   X   V       W   G   L    ����                                                                                                                                                                                                                                                                                                                            G   L       G   V       v   V    ^1     �   F   H   `      Z                        m_axis_tdata_tb  <= std_logic_vector(to_signed(data,data'length));5�_�   W   Y           X   >        ����                                                                                                                                                                                                                                                                                                                            >   V       >   V       V   V    ^;     �   =   ?   _    �   >   ?   _    �   =   >          W                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,data'length));5�_�   X   Z           Y   >       ����                                                                                                                                                                                                                                                                                                                            >           >   d       V   V    ^=   	 �   =   ?          e                        m_axis_tdata_tb  <= std_logic_vector(to_signed(data,m_axis_tdata_tb'length));5�_�   Y   [           Z   !   <    ����                                                                                                                                                                                                                                                                                                                            !   <       !   E       v   E    ^�     �       "   `      G   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):="01110111";5�_�   Z   \           [   !   <    ����                                                                                                                                                                                                                                                                                                                            !   <       !   E       v   E    ^�     �       "   `      J   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');5�_�   [   ]           \   >   I    ����                                                                                                                                                                                                                                                                                                                            >   I       >   ^       v   ^    ^�     �   =   ?   `      b                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,m_axis_tdata_tb'length));5�_�   \   ^           ]   G        ����                                                                                                                                                                                                                                                                                                                            G   I       G   I       V   I    ^�     �   F   H   _    �   G   H   _    �   F   G          e                        m_axis_tdata_tb  <= std_logic_vector(to_signed(data,m_axis_tdata_tb'length));5�_�   ]   _           ^   G       ����                                                                                                                                                                                                                                                                                                                            G           G   L       V   I    ^�   
 �   F   H          M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   ^   `           _   >   )    ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   =   ?   `      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   _   a           `   G       ����                                                                                                                                                                                                                                                                                                                                                             ^�     �   F   H   `    �   G   H   `    5�_�   `   b           a   H       ����                                                                                                                                                                                                                                                                                                                                                             ^�    �   G   I   a      P                        m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   a   c           b   Z       ����                                                                                                                                                                                                                                                                                                                            Z          ]                 ^	(     �   Y   ^   a      -           s_axis_tdata  =>s_axis_tdata_tb  ,   -           s_axis_tvalid =>s_axis_tvalid_tb ,   -           s_axis_tlast  =>s_axis_tlast_tb  ,   -           s_axis_tready =>s_axis_tready_tb ,5�_�   b   d           c   V       ����                                                                                                                                                                                                                                                                                                                            V          Y                 ^	,    �   U   Z   a      -           m_axis_tdata  =>m_axis_tdata_tb  ,   -           m_axis_tvalid =>m_axis_tvalid_tb ,   -           m_axis_tlast  =>m_axis_tlast_tb  ,   -           m_axis_tready =>m_axis_tready_tb ,5�_�   c   e           d   %        ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	     �   $   )   a    �   %   &   a    5�_�   d   f           e   %       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   $   &   e      K   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   e   g           f   &       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   %   '   e      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';5�_�   f   h           g   '       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   &   (   e      ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';5�_�   g   i           h   (       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   '   )   e      ,   signal s_axis_tready_tb : STD_LOGIC:='0';5�_�   h   j           i   (   ,    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   '   )   e      /   signal s_axis_tready_empty : STD_LOGIC:='0';5�_�   i   k           j   &   ,    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   %   '   e      /   signal s_axis_tvalid_empty : STD_LOGIC:='1';5�_�   j   l           k   Z   (    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   Y   [   e      -           m_axis_tdata  =>s_axis_tdata_tb  ,5�_�   k   m           l   [   )    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   Z   \   e      -           m_axis_tvalid =>s_axis_tvalid_tb ,5�_�   l   n           m   \   (    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�     �   [   ]   e      -           m_axis_tlast  =>s_axis_tlast_tb  ,5�_�   m   o           n   ]   )    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�    �   \   ^   e      -           m_axis_tready =>s_axis_tready_tb ,5�_�   n   p           o   $       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^	�    �   $   &   e    5�_�   o   q           p   D       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
:    �   C   E   f      2                     data             := data + 1;5�_�   p   r           q   D       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
S     �   C   E   f      4                     --data             := data + 1;5�_�   q   s           r   D       ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
S     �   C   E   f      3                     -data             := data + 1;5�_�   r   t           s   3   #    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
`     �   2   4   f      2      variable data :integer range -128 to 127:=0;5�_�   s   u           t   3   (    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
d    �   2   4   f      /      variable data :integer range 0 to 127:=0;5�_�   t   v           u   D   )    ����                                                                                                                                                                                                                                                                                                                            !          $          V       ^
�     �   C   E   f      2                     data             := data + 1;5�_�   u   w           v   D   (    ����                                                                                                                                                                                                                                                                                                                            D   (       D   3       v   3    ^
�     �   C   E   f      =                     data             := to_integer(data + 1;5�_�   v   x           w   3   #    ����                                                                                                                                                                                                                                                                                                                            3   #       3   *       v   *    ^
�     �   2   4   f      /      variable data :integer range 0 to 255:=0;5�_�   w   y           x   3   #    ����                                                                                                                                                                                                                                                                                                                            3   #       3   *       v   *    ^
�    �   2   4   f      '      variable data :integer range :=0;5�_�   x   z           y   3       ����                                                                                                                                                                                                                                                                                                                            3          3   $       v   $    ^
�    �   2   4   f      )      variable data :integer range <>:=0;5�_�   y   {           z   C   )    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^
�    �   B   D   f      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));5�_�   z   |           {   D   (    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^
�     �   C   E   f      1                     data             :=data + 1;5�_�   {   }           |   D   ;    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^
�    �   C   E   f      <                     data             :=to_integer(data + 1;5�_�   |   ~           }   D   ;    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^
�     �   C   E   f      ?                     data             :=to_integer(data + 1,8);5�_�   }   �           ~   D   ;    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^
�    �   C   E   f      >                     data             :=to_integer(data + 18);5�_�   ~   �          �   3       ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^3     �   2   4   f             variable data :integer:=0;5�_�   �   �           �   D   +    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^R     �   C   E   f      =                     data             :=to_integer(data + 1);5�_�   �   �           �   D   :    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^U     �   C   E   f      <                     data             :=to_signed(data + 1);5�_�   �   �           �   D   (    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^`     �   C   E   f      >                     data             :=to_signed(data + 1,8);5�_�   �   �           �   D   H    ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^d    �   C   E   f      I                     data             :=to_integer(to_signed(data + 1,8);5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^�    �   ]   _          0           m_axis_tready =>s_axis_tready_empty ,�   \   ^          0           m_axis_tlast  =>s_axis_tlast_empty  ,�   [   ]          0           m_axis_tvalid =>s_axis_tvalid_empty ,�   Z   \          0           m_axis_tdata  =>s_axis_tdata_empty  ,�   (   *          /   signal s_axis_tready_empty : STD_LOGIC:='1';�   '   )          /   signal s_axis_tlast_empty  : STD_LOGIC:='0';�   &   (          /   signal s_axis_tvalid_empty : STD_LOGIC:='0';�   %   '          N   signal s_axis_tdata_empty  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �   �           �            ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^     �                  5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       #                 ^     �       $   e      ,   signal s_axis_tvalid_tb : STD_LOGIC:='1';   ,   signal s_axis_tlast_tb  : STD_LOGIC:='0';   ,   signal s_axis_tready_tb : STD_LOGIC:='0';�      !   e      K   signal s_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                       ^#     �          e      ,   signal m_axis_tvalid_tb : STD_LOGIC:='0';   ,   signal m_axis_tlast_tb  : STD_LOGIC:='0';   ,   signal m_axis_tready_tb : STD_LOGIC:='1';�         e      J   signal m_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       #                 ^O     �      $   e      L   signal si_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');   -   signal si_axis_tvalid_tb : STD_LOGIC:='1';   -   signal si_axis_tlast_tb  : STD_LOGIC:='0';   -   signal si_axis_tready_tb : STD_LOGIC:='0';5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            ^          a                 ^^     �   ^   b   e      -           s_axis_tvalid =>m_axis_tvalid_tb ,   -           s_axis_tlast  =>m_axis_tlast_tb  ,   -           s_axis_tready =>m_axis_tready_tb ,�   ]   _   e      -           s_axis_tdata  =>m_axis_tdata_tb  ,5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^d     �   Z   ^   e      1           m_axis_tvalid =>s_axis_tvalid_output ,   1           m_axis_tlast  =>s_axis_tlast_output  ,   1           m_axis_tready =>s_axis_tready_output ,�   Y   [   e      1           m_axis_tdata  =>s_axis_tdata_output  ,5�_�   �   �           �   Z   (    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^h     �   Y   [   e      2           m_axis_tdata  =>s2_axis_tdata_output  ,5�_�   �   �           �   [   )    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^i     �   Z   \   e      2           m_axis_tvalid =>s2_axis_tvalid_output ,5�_�   �   �           �   \   (    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^j     �   [   ]   e      2           m_axis_tlast  =>s2_axis_tlast_output  ,5�_�   �   �           �   ]   )    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^k     �   \   ^   e      2           m_axis_tready =>s2_axis_tready_output ,5�_�   �   �           �   ^   (    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^l     �   ]   _   e      .           s_axis_tdata  =>m1_axis_tdata_tb  ,5�_�   �   �           �   _   )    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^m     �   ^   `   e      .           s_axis_tvalid =>m1_axis_tvalid_tb ,5�_�   �   �   �       �   `   (    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^p     �   _   a   e      .           s_axis_tlast  =>m1_axis_tlast_tb  ,5�_�   �   �           �   a   )    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^p     �   `   b   e      .           s_axis_tready =>m1_axis_tready_tb ,5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^{     �   %   )   e      0   signal s_axis_tvalid_output : STD_LOGIC:='0';   0   signal s_axis_tlast_output  : STD_LOGIC:='0';   0   signal s_axis_tready_output : STD_LOGIC:='1';�   $   &   e      O   signal s_axis_tdata_output  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^}     �   $   &   e      P   signal s2_axis_tdata_output  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^~     �   %   '   e      1   signal s2_axis_tvalid_output : STD_LOGIC:='0';5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^~     �   &   (   e      1   signal s2_axis_tlast_output  : STD_LOGIC:='0';5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^     �   '   )   e      1   signal s2_axis_tready_output : STD_LOGIC:='1';5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            %          *          V       ^�     �   b   d   e      .           rst           =>rst_tb           );�   a   c   e      -           clk           =>clk_tb           ,�   `   b   e      *           s_axis_tready =>m1_axis_tready,�   _   a   e      )           s_axis_tlast  =>m1_axis_tlast,�   ^   `   e      *           s_axis_tvalid =>m1_axis_tvalid,�   ]   _   e      )           s_axis_tdata  =>m1_axis_tdata,�   \   ^   e      *           m_axis_tready =>s2_axis_tready,�   [   ]   e      )           m_axis_tlast  =>s2_axis_tlast,�   Z   \   e      *           m_axis_tvalid =>s2_axis_tvalid,�   Y   [   e      )           m_axis_tdata  =>s2_axis_tdata,�   X   Z   e          port map(  �   U   W   e         end process axi_master_proc;�   T   V   e            end if;�   S   U   e               end if;�   R   T   e                  end case;�   Q   S   e                        end if;�   P   R   e                           end if;�   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   N   P   e      0                        s_axis_tready_tb <= '1';�   M   O   e      0                        m_axis_tvalid_tb <= '0';�   L   N   e                           else�   K   M   e      R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   J   L   e      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));�   I   K   e      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   H   J   e      Q                     bitCounter := bitCounter+1;                     --incremento�   G   I   e      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   F   H   e      $               when waitingMready =>�   E   G   e                        end if;�   D   F   e      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   C   E   e      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   B   D   e      J                     data             :=to_integer(to_signed(data + 1,8));�   A   C   e      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   @   B   e      +                     bitCounter       := 0;�   ?   A   e      -                     s_axis_tready_tb <= '0';�   >   @   e      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   =   ?   e      $               when waitingSvalid =>�   <   >   e                  case state is�   ;   =   e               else�   :   <   e                  data  := 0;�   9   ;   e      0            m_axis_tdata_tb  <= (others => '0');�   8   :   e      $            m_axis_tvalid_tb <= '0';�   7   9   e      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato�   6   8   e      $            s_axis_tready_tb <= '1';�   5   7   e      +            state         <= waitingSvalid;�   4   6   e               if rst_tb = '0' then�   3   5   e      !      if rising_edge(clk_tb) then�   2   4   e         begin�   1   3   e      2      variable data :integer range -128 to 127:=0;�   0   2   e      0      variable bitCounter :integer range 0 to 8;�   /   1   e      &   axi_master_proc:process (clk_tb) is�   -   /   e          rst_tb   <= '1' after 180 ns;�   ,   .   e      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   )   +   e      :   signal rst_tb          :                STD_LOGIC:='0';�   (   *   e      :   signal clk_tb          :                STD_LOGIC:='0';�   '   )   e      )   signal s2_axis_tready: STD_LOGIC:='1';�   &   (   e      )   signal s2_axis_tlast:  STD_LOGIC:='0';�   %   '   e      )   signal s2_axis_tvalid: STD_LOGIC:='0';�   $   &   e      H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   "   $   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�   !   #   e      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';�       "   e      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';�      !   e      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�          e      -   signal m1_axis_tready_tb : STD_LOGIC:='1';�         e      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';�         e      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';�         e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         e         end component split_1to8;�         e      *           rst           : in  STD_LOGIC);�         e      )           clk           : in  STD_LOGIC;�         e      )           s_axis_tready : out STD_LOGIC;�         e      )           s_axis_tlast  : in  STD_LOGIC;�         e      )           s_axis_tvalid : in  STD_LOGIC;�         e      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         e      )           m_axis_tready : in  STD_LOGIC;�         e      )           m_axis_tlast  : out STD_LOGIC;�         e      )           m_axis_tvalid : out STD_LOGIC;�         e      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         e      	    port(�         e         component split_1to8 is�   	      e      +   signal state:axiStates := waitingSvalid;�      
   e      4   type axiStates is (waitingSvalid, waitingMready);�   )   +          ,   signal rst_tb           : STD_LOGIC:='0';�   &   (          (   signal s2_axis_tlast: STD_LOGIC:='0';�   %   '          )   signal s2_axis_tvalid: STD_LOGIC:='0';�   $   &          G   signal s2_axis_tdata: STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   (   *          ,   signal clk_tb           : STD_LOGIC:='0';�   '   )          )   signal s2_axis_tready: STD_LOGIC:='1';5�_�   �   �   �       �   '        ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   &   (          )   signal s2_axis_tlast:  STD_LOGIC:='0';�   %   '          )   signal s2_axis_tvalid: STD_LOGIC:='0';�   $   &          H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   $   &   e      I   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   &   (   e      >   signal s2_axis_tlast:  STD_LOGIC:                     ='0';5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   &   (   e      ?   signal s2_axis_tlast :  STD_LOGIC:                     ='0';5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   &   (   e      @   signal s2_axis_tlast :i  STD_LOGIC:                     ='0';5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                            %          (                 ^�     �   %   )   e      >   signal s2_axis_tvalid: STD_LOGIC:                     ='0';   ?   signal s2_axis_tlast :  STD_LOGIC:                     ='0';   )   signal s2_axis_tready: STD_LOGIC:='1';�   $   &   e      J   signal s2_axis_tdata :  STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            )          *                 ^�     �   )   +   e      :   signal rst_tb          :                STD_LOGIC:='0';�   (   *   e      :   signal clk_tb          :                STD_LOGIC:='0';5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                            %          *          V       ^�     �   b   d   e      .           rst           =>rst_tb           );�   a   c   e      -           clk           =>clk_tb           ,�   `   b   e      *           s_axis_tready =>m1_axis_tready,�   _   a   e      )           s_axis_tlast  =>m1_axis_tlast,�   ^   `   e      *           s_axis_tvalid =>m1_axis_tvalid,�   ]   _   e      )           s_axis_tdata  =>m1_axis_tdata,�   \   ^   e      *           m_axis_tready =>s2_axis_tready,�   [   ]   e      )           m_axis_tlast  =>s2_axis_tlast,�   Z   \   e      *           m_axis_tvalid =>s2_axis_tvalid,�   Y   [   e      )           m_axis_tdata  =>s2_axis_tdata,�   X   Z   e          port map(  �   U   W   e         end process axi_master_proc;�   T   V   e            end if;�   S   U   e               end if;�   R   T   e                  end case;�   Q   S   e                        end if;�   P   R   e                           end if;�   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   N   P   e      0                        s_axis_tready_tb <= '1';�   M   O   e      0                        m_axis_tvalid_tb <= '0';�   L   N   e                           else�   K   M   e      R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   J   L   e      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));�   I   K   e      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   H   J   e      Q                     bitCounter := bitCounter+1;                     --incremento�   G   I   e      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   F   H   e      $               when waitingMready =>�   E   G   e                        end if;�   D   F   e      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   C   E   e      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   B   D   e      J                     data             :=to_integer(to_signed(data + 1,8));�   A   C   e      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   @   B   e      +                     bitCounter       := 0;�   ?   A   e      -                     s_axis_tready_tb <= '0';�   >   @   e      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   =   ?   e      $               when waitingSvalid =>�   <   >   e                  case state is�   ;   =   e               else�   :   <   e                  data  := 0;�   9   ;   e      0            m_axis_tdata_tb  <= (others => '0');�   8   :   e      $            m_axis_tvalid_tb <= '0';�   7   9   e      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato�   6   8   e      $            s_axis_tready_tb <= '1';�   5   7   e      +            state         <= waitingSvalid;�   4   6   e               if rst_tb = '0' then�   3   5   e      !      if rising_edge(clk_tb) then�   2   4   e         begin�   1   3   e      2      variable data :integer range -128 to 127:=0;�   0   2   e      0      variable bitCounter :integer range 0 to 8;�   /   1   e      &   axi_master_proc:process (clk_tb) is�   -   /   e          rst_tb   <= '1' after 180 ns;�   ,   .   e      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   )   +   e      *   signal rst_tb         : STD_LOGIC:='0';�   (   *   e      *   signal clk_tb         : STD_LOGIC:='0';�   '   )   e      *   signal s2_axis_tready : STD_LOGIC:='1';�   &   (   e      1   signal s2_axis_tlast  : STD_LOGIC:       ='0';�   %   '   e      1   signal s2_axis_tvalid : STD_LOGIC:       ='0';�   $   &   e      J   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');�   "   $   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�   !   #   e      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';�       "   e      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';�      !   e      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�          e      -   signal m1_axis_tready_tb : STD_LOGIC:='1';�         e      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';�         e      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';�         e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         e         end component split_1to8;�         e      *           rst           : in  STD_LOGIC);�         e      )           clk           : in  STD_LOGIC;�         e      )           s_axis_tready : out STD_LOGIC;�         e      )           s_axis_tlast  : in  STD_LOGIC;�         e      )           s_axis_tvalid : in  STD_LOGIC;�         e      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         e      )           m_axis_tready : in  STD_LOGIC;�         e      )           m_axis_tlast  : out STD_LOGIC;�         e      )           m_axis_tvalid : out STD_LOGIC;�         e      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         e      	    port(�         e         component split_1to8 is�   	      e      +   signal state:axiStates := waitingSvalid;�      
   e      4   type axiStates is (waitingSvalid, waitingMready);�   )   +          ;   signal rst_tb           :                STD_LOGIC:='0';�   &   (          B   signal s2_axis_tlast    :  STD_LOGIC:                     ='0';�   %   '          A   signal s2_axis_tvalid   : STD_LOGIC:                     ='0';�   $   &          M   signal s2_axis_tdata    :  STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');�   (   *          ;   signal clk_tb           :                STD_LOGIC:='0';�   '   )          ,   signal s2_axis_tready   : STD_LOGIC:='1';5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                            &   %       *   %       V   %    ^�     �   b   d   e      .           rst           =>rst_tb           );�   a   c   e      -           clk           =>clk_tb           ,�   `   b   e      *           s_axis_tready =>m1_axis_tready,�   _   a   e      )           s_axis_tlast  =>m1_axis_tlast,�   ^   `   e      *           s_axis_tvalid =>m1_axis_tvalid,�   ]   _   e      )           s_axis_tdata  =>m1_axis_tdata,�   \   ^   e      *           m_axis_tready =>s2_axis_tready,�   [   ]   e      )           m_axis_tlast  =>s2_axis_tlast,�   Z   \   e      *           m_axis_tvalid =>s2_axis_tvalid,�   Y   [   e      )           m_axis_tdata  =>s2_axis_tdata,�   X   Z   e          port map(  �   U   W   e         end process axi_master_proc;�   T   V   e            end if;�   S   U   e               end if;�   R   T   e                  end case;�   Q   S   e                        end if;�   P   R   e                           end if;�   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   N   P   e      0                        s_axis_tready_tb <= '1';�   M   O   e      0                        m_axis_tvalid_tb <= '0';�   L   N   e                           else�   K   M   e      R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   J   L   e      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));�   I   K   e      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   H   J   e      Q                     bitCounter := bitCounter+1;                     --incremento�   G   I   e      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   F   H   e      $               when waitingMready =>�   E   G   e                        end if;�   D   F   e      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   C   E   e      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   B   D   e      J                     data             :=to_integer(to_signed(data + 1,8));�   A   C   e      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   @   B   e      +                     bitCounter       := 0;�   ?   A   e      -                     s_axis_tready_tb <= '0';�   >   @   e      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   =   ?   e      $               when waitingSvalid =>�   <   >   e                  case state is�   ;   =   e               else�   :   <   e                  data  := 0;�   9   ;   e      0            m_axis_tdata_tb  <= (others => '0');�   8   :   e      $            m_axis_tvalid_tb <= '0';�   7   9   e      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato�   6   8   e      $            s_axis_tready_tb <= '1';�   5   7   e      +            state         <= waitingSvalid;�   4   6   e               if rst_tb = '0' then�   3   5   e      !      if rising_edge(clk_tb) then�   2   4   e         begin�   1   3   e      2      variable data :integer range -128 to 127:=0;�   0   2   e      0      variable bitCounter :integer range 0 to 8;�   /   1   e      &   axi_master_proc:process (clk_tb) is�   -   /   e          rst_tb   <= '1' after 180 ns;�   ,   .   e      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   )   +   e      -   signal rst_tb         : STD_LOGIC  := '0';�   (   *   e      -   signal clk_tb         : STD_LOGIC  := '0';�   '   )   e      -   signal s2_axis_tready : STD_LOGIC  := '1';�   &   (   e      -   signal s2_axis_tlast  : STD_LOGIC:  = '0';�   %   '   e      -   signal s2_axis_tvalid : STD_LOGIC:  = '0';�   $   &   e      J   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');�   "   $   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�   !   #   e      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';�       "   e      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';�      !   e      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�          e      -   signal m1_axis_tready_tb : STD_LOGIC:='1';�         e      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';�         e      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';�         e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         e         end component split_1to8;�         e      *           rst           : in  STD_LOGIC);�         e      )           clk           : in  STD_LOGIC;�         e      )           s_axis_tready : out STD_LOGIC;�         e      )           s_axis_tlast  : in  STD_LOGIC;�         e      )           s_axis_tvalid : in  STD_LOGIC;�         e      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         e      )           m_axis_tready : in  STD_LOGIC;�         e      )           m_axis_tlast  : out STD_LOGIC;�         e      )           m_axis_tvalid : out STD_LOGIC;�         e      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         e      	    port(�         e         component split_1to8 is�   	      e      +   signal state:axiStates := waitingSvalid;�      
   e      4   type axiStates is (waitingSvalid, waitingMready);�   %   '          1   signal s2_axis_tvalid : STD_LOGIC:       ='0';�   &   (          1   signal s2_axis_tlast  : STD_LOGIC:       ='0';�   )   +          *   signal rst_tb         : STD_LOGIC:='0';�   (   *          *   signal clk_tb         : STD_LOGIC:='0';�   '   )          *   signal s2_axis_tready : STD_LOGIC:='1';5�_�   �   �           �   &   $    ����                                                                                                                                                                                                                                                                                                                            &   $       '   $          $    ^�     �   &   (   e      -   signal s2_axis_tlast  : STD_LOGIC:  = '0';�   %   '   e      -   signal s2_axis_tvalid : STD_LOGIC:  = '0';5�_�   �   �           �   &   &    ����                                                                                                                                                                                                                                                                                                                            &   &       '   '          '    ^�     �   %   (   e      1   signal s2_axis_tvalid : STD_LOGIC   l:  = '0';   1   signal s2_axis_tlast  : STD_LOGIC   l:  = '0';5�_�   �   �           �   &   '    ����                                                                                                                                                                                                                                                                                                                            &   '       '   (          (    ^�     �   %   (   e      /   signal s2_axis_tvalid : STD_LOGIC  :  = '0';   /   signal s2_axis_tlast  : STD_LOGIC  :  = '0';5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            )          *          V       ^�     �   (   )          -   signal clk_tb         : STD_LOGIC  := '0';   -   signal rst_tb         : STD_LOGIC  := '0';5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�     �         c    �         c    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      -   signal rst_tb         : STD_LOGIC  := '0';�         e      -   signal clk_tb         : STD_LOGIC  := '0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      /   signal rst_tb           : STD_LOGIC  := '0';�         e      /   signal clk_tb           : STD_LOGIC  := '0';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      0   signal rst_tb            : STD_LOGIC  := '0';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      0   signal clk_tb            : STD_LOGIC  := '0';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      /   signal rst_tb            : STD_LOGIC := '0';5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e      /   signal clk_tb            : STD_LOGIC := '0';5�_�   �   �   �       �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e    5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            8          ;                 ^     �   8   <   f      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato   $            m_axis_tvalid_tb <= '0';   0            m_axis_tdata_tb  <= (others => '0');�   7   9   f      $            s_axis_tready_tb <= '1';5�_�   �   �           �   8       ����                                                                                                                                                                                                                                                                                                                            8          ;                 ^	     �   7   9   f      %            s1_axis_tready_tb <= '1';5�_�   �   �           �   9       ����                                                                                                                                                                                                                                                                                                                            8          ;                 ^	     �   8   :   f      U            s1_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   �   �           �   :       ����                                                                                                                                                                                                                                                                                                                            8          ;                 ^
     �   9   ;   f      %            m1_axis_tvalid_tb <= '0';5�_�   �   �           �   ;       ����                                                                                                                                                                                                                                                                                                                            8          ;                 ^
     �   :   <   f      1            m1_axis_tdata_tb  <= (others => '0');5�_�   �   �           �   @       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   @   B   f      -                     s_axis_tready_tb <= '0';�   ?   A   f      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo5�_�   �   �           �   @   #    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   ?   A   f      v                  if s1_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo5�_�   �   �           �   A   #    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   @   B   f      .                     s1_axis_tready_tb <= '0';5�_�   �   �           �   C       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   B   D   f      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   �   �           �   C   "    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   B   D   f      N                     m1_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   �   �           �   E       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   D   F   f      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   �   �           �   E   #    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^     �   D   F   f      s                     m1_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^!     �   H   J   f      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�   �   �           �   I   #    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^#     �   H   J   f      u                  if m1_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^&     �   K   M   f      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            @          A                 ^(     �   K   M   f      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));5�_�   �   �           �   L   "    ����                                                                                                                                                                                                                                                                                                                            @          A                 ^*     �   K   M   f      [                     m1_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));5�_�   �   �           �   L   %    ����                                                                                                                                                                                                                                                                                                                            L   %       L   1       v   1    ^<     �   K   M   f      V                     m1_axis_tdata<= "10101111";--std_logic_vector(to_signed(data,8));5�_�   �   �           �   L        ����                                                                                                                                                                                                                                                                                                                            L   %       L   %       V   %    ^B     �   K   M   e    �   L   M   e    �   K   L          I                     m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            L           L   H       V   %    ^D     �   L   M          R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            L           L   H       V   %    ^D     �   K   M          I                     m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            O          N                 ^I     �   N   P   e      0                        s_axis_tready_tb <= '1';�   M   O   e      0                        m_axis_tvalid_tb <= '0';5�_�   �   �           �   N   &    ����                                                                                                                                                                                                                                                                                                                            N   &       O   (          (    ^L     �   M   P   e      1                        m1_axis_tvalid_tb <= '0';   1                        s1_axis_tready_tb <= '1';5�_�   �   �           �   P   &    ����                                                                                                                                                                                                                                                                                                                            N   &       O   (          (    ^M     �   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �   P   &    ����                                                                                                                                                                                                                                                                                                                            N   &       O   (          (    ^M     �   O   Q   e      �                        state           <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                  V        ^]     �         e         end component split_1to8;�         e         component split_1to8 is5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       &           V        ^b     �   %   '   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�          e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                            (           +           V        ^e     �   *   ,   e      -   signal s2_axis_tready : STD_LOGIC  := '1';�   '   )   e      J   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                            (           +           V        ^f     �   &   '           5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            '           *           V        ^g     �                 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            &           )           V        ^h     �                 5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                            %           (           V        ^m     �      
   b      4   type axiStates is (waitingSvalid, waitingMready);5�_�   �   �           �   
       ����                                                                                                                                                                                                                                                                                                                            %           (           V        ^o     �   	      b      +   signal state:axiStates := waitingSvalid;5�_�   �   �           �   U        ����                                                                                                                                                                                                                                                                                                                            U          `          V       ^y    �   _   a   b      .           rst           =>rst_tb           );�   T   V   b      split_1to8_inst:split_1to85�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            U          `          V       ^�     �         b      !   component split_1to8 is/*{{{*/5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            U          `          V       ^�    �         b      #   end component split_1to8;/*}}}*/5�_�   �   �           �      K    ����                                                                                                                                                                                                                                                                                                                            U          `          V       ^�     �         b      N   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�   �   �           �   $   -    ����                                                                                                                                                                                                                                                                                                                            U          `          V       ^�     �   #   %   b      4   signal s1_axis_tready_tb : STD_LOGIC:='0';/*}}}*/5�_�   �   �           �      ,    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�         b      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');5�_�   �   �           �      K    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      N   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�   �   �           �   $   2    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      4   signal s1_axis_tready_tb : STD_LOGIC:='0';/*}}}*/5�_�   �   �           �   $   2    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      3   signal s1_axis_tready_tb : STD_LOGIC:='0';/*}}}/5�_�   �   �           �   $   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      2   signal s1_axis_tready_tb : STD_LOGIC:='0';/*}}}5�_�   �   �           �   $   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      1   signal s1_axis_tready_tb : STD_LOGIC:='0';*}}}5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      &   end component split_1to8; --/*}}}*/5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      %   end component split_1to8; --*}}}*/5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      $   end component split_1to8; --}}}*/5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      #   end component split_1to8; --}}}/5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      $   component split_1to8 is --/*{{{*/5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      #   component split_1to8 is --*{{{*/5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �         b      "   component split_1to8 is --{{{*/5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�    �         b      !   component split_1to8 is --{{{/5�_�   �   �           �   $   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   #   %   b      0   signal s1_axis_tready_tb : STD_LOGIC:='0';}}}5�_�   �   �           �   $   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�    �   #   %   b      2   signal s1_axis_tready_tb : STD_LOGIC:='0';--}}}5�_�   �   �           �   %   J    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   $   &   b      M   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');{{{5�_�   �   �           �   (   3    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   '   )   b      4   signal s2_axis_tready : STD_LOGIC  := '1';/*}}}*/5�_�   �   �           �   (   2    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   '   )   b      3   signal s2_axis_tready : STD_LOGIC  := '1';/*}}}*5�_�   �   �           �   (   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   '   )   b      2   signal s2_axis_tready : STD_LOGIC  := '1';/*}}}5�_�   �   �           �   (   -    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�    �   '   )   b      2   signal s2_axis_tready : STD_LOGIC  := '1';--}}}5�_�   �   �           �   %   J    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   $   '   b      P   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0'); --{{{5�_�   �   �           �   %   8    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   $   &   c      J   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');5�_�   �   �           �   %   :    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   $   &   c      K   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0) : = (others=>'0');5�_�   �   �           �   %   :    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�   ! �   $   &   c      J   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0) := (others=>'0');      --{{{5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   T   V   b      !split_1to8_inst:split_1to8/*{{{*/5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   T   V   b      $split_1to8_inst:split_1to8 --/*{{{*/5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   T   V   b      #split_1to8_inst:split_1to8 --*{{{*/5�_�   �   �           �   U        ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   T   V   b      "split_1to8_inst:split_1to8 --{{{*/5�_�   �   �           �   U        ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^�     �   T   V   b      !split_1to8_inst:split_1to8 --{{{/5�_�   �   �           �   `   .    ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^   " �   _   a   b      1           rst           =>rst_tb           );}}}5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �         b      Q   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �         b      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �          b      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �      !   b      -   signal m1_axis_tready_tb : STD_LOGIC:='1';5�_�   �              �   !       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �       "   b      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�   �                "       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �   !   #   b      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';5�_�                  #       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �   "   $   b      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';5�_�                 $       ����                                                                                                                                                                                                                                                                                                                            $   ,          ,       V   ,    ^     �   #   %   b      3   signal s1_axis_tready_tb : STD_LOGIC:='0'; --}}}5�_�                         ����                                                                                                                                                                                                                                                                                                                            $                    V       ^   $ �   _   a   b      4           rst           =>rst_tb           ); --}}}�   ^   `   b      -           clk           =>clk_tb           ,�   ]   _   b      *           s_axis_tready =>m1_axis_tready,�   \   ^   b      )           s_axis_tlast  =>m1_axis_tlast,�   [   ]   b      *           s_axis_tvalid =>m1_axis_tvalid,�   Z   \   b      )           s_axis_tdata  =>m1_axis_tdata,�   Y   [   b      *           m_axis_tready =>s2_axis_tready,�   X   Z   b      )           m_axis_tlast  =>s2_axis_tlast,�   W   Y   b      *           m_axis_tvalid =>s2_axis_tvalid,�   V   X   b      )           m_axis_tdata  =>s2_axis_tdata,�   U   W   b          port map(  �   R   T   b         end process axi_master_proc;�   Q   S   b            end if;�   P   R   b               end if;�   O   Q   b                  end case;�   N   P   b                        end if;�   M   O   b                           end if;�   L   N   b      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   K   M   b      .                        s1_axis_tready <= '1';�   J   L   b      .                        m1_axis_tvalid <= '0';�   I   K   b                           else�   H   J   b      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   G   I   b      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   F   H   b      Q                     bitCounter := bitCounter+1;                     --incremento�   E   G   b      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   D   F   b      $               when waitingMready =>�   C   E   b                        end if;�   B   D   b      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   A   C   b      o                     m1_axis_tvalid<= '1';                         --como puedo mandar, le avoso que tengo dato�   @   B   b      J                     data             :=to_integer(to_signed(data + 1,8));�   ?   A   b      I                     m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   >   @   b      +                     bitCounter       := 0;�   =   ?   b      *                     s1_axis_tready<= '0';�   <   >   b      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   ;   =   b      $               when waitingSvalid =>�   :   <   b                  case state is�   9   ;   b               else�   8   :   b                  data  := 0;�   7   9   b      ,            m1_axis_tdata<= (others => '0');�   6   8   b      !            m1_axis_tvalid<= '0';�   5   7   b      Q            s1_axis_tvalid<= '1'; --que haga de cuentqa que siempre tiene un dato�   4   6   b      !            s1_axis_tready<= '1';�   3   5   b      +            state         <= waitingSvalid;�   2   4   b               if rst_tb = '0' then�   1   3   b      !      if rising_edge(clk_tb) then�   0   2   b         begin�   /   1   b      2      variable data :integer range -128 to 127:=0;�   .   0   b      0      variable bitCounter :integer range 0 to 8;�   -   /   b      &   axi_master_proc:process (clk_tb) is�   +   -   b          rst_tb   <= '1' after 180 ns;�   *   ,   b      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   '   )   b      3   signal s2_axis_tready : STD_LOGIC  := '1'; --}}}�   &   (   b      -   signal s2_axis_tlast  : STD_LOGIC  := '0';�   %   '   b      -   signal s2_axis_tvalid : STD_LOGIC  := '0';�   $   &   b      P   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0) := (others=>'0'); --{{{�   #   %   b      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   "   $   b      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   !   #   b      )   signal s1_axis_tvalid: STD_LOGIC:='1';�       "   b      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�      !   b      )   signal m1_axis_tready: STD_LOGIC:='1';�          b      )   signal m1_axis_tlast:  STD_LOGIC:='0';�         b      )   signal m1_axis_tvalid: STD_LOGIC:='0';�         b      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�         b      .   signal rst_tb            : STD_LOGIC:= '0';�         b      .   signal clk_tb            : STD_LOGIC:= '0';�         b      "   end component split_1to8; --}}}�         b      *           rst           : in  STD_LOGIC);�         b      )           clk           : in  STD_LOGIC;�         b      )           s_axis_tready : out STD_LOGIC;�         b      )           s_axis_tlast  : in  STD_LOGIC;�         b      )           s_axis_tvalid : in  STD_LOGIC;�         b      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         b      )           m_axis_tready : in  STD_LOGIC;�         b      )           m_axis_tlast  : out STD_LOGIC;�         b      )           m_axis_tvalid : out STD_LOGIC;�         b      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         b      	    port(�         b          component split_1to8 is --{{{�   	      b      .   signal state   :axiStates := waitingSvalid;�      
   b      6   type   axiStates is (waitingSvalid, waitingMready);�                )   signal m1_axis_tvalid: STD_LOGIC:='0';�   !   #          )   signal s1_axis_tvalid: STD_LOGIC:='1';�   #   %          /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   "   $          (   signal s1_axis_tlast: STD_LOGIC:='0';�                L   signal m1_axis_tdata: STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�       "          G   signal s1_axis_tdata: STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�      !          )   signal m1_axis_tready: STD_LOGIC:='1';�                 (   signal m1_axis_tlast: STD_LOGIC:='0';5�_�                 .        ����                                                                                                                                                                                                                                                                                                                            .           S           V        ^7     �   R   T   b         end process axi_master_proc;�   -   /   b      &   axi_master_proc:process (clk_tb) is5�_�                 T        ����                                                                                                                                                                                                                                                                                                                            .           S           V        ^8     �   S   T           5�_�                         ����                                                                                                                                                                                                                                                                                                                            .           S           V        ^C     �         a    �         a    5�_�                         ����                                                                                                                                                                                                                                                                                                                                       )   "       V        ^e     �   (   *          "   end component split_1to8; --}}}�                    component split_1to8 is --{{{5�_�    	             c        ����                                                                                                                                                                                                                                                                                                                                       )   "       V        ^l     �   b   o   p    �   c   d   p    5�_�    
          	   o        ����                                                                                                                                                                                                                                                                                                                            o           z   4       V        ^n     �   n   p           split_1to8_inst:split_1to8 --{{{5�_�  	            
   b       ����                                                                                                                                                                                                                                                                                                                            o           z   4       V        ^x     �   b   d   |    5�_�  
               <        ����                                                                                                                                                                                                                                                                                                                            p           {   4       V        ^y     �   ;   <           5�_�                         ����                                                                                                                                                                                                                                                                                                                            o           z   4       V        ^�     �                 5�_�                         ����                                                                                                                                                                                                                                                                                                                            n           y   4       V        ^�     �                 5�_�                         ����                                                                                                                                                                                                                                                                                                                            m           x   4       V        ^�     �         {       �         z    5�_�                         ����                                                                                                                                                                                                                                                                                                                            n           y   4       V        ^�     �         {    5�_�                         ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         |      end;�          |      library ieee;5�_�                 ,        ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �   +   4   |    �   ,   -   |    5�_�                 4        ����                                                                                                                                                                                                                                                                                                                            4           ;   /       V        ^�     �   6   8          )   signal m1_axis_tready: STD_LOGIC:='1';�   5   7          )   signal m1_axis_tlast:  STD_LOGIC:='0';�   4   6          )   signal m1_axis_tvalid: STD_LOGIC:='0';�   3   5          M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�                 8        ����                                                                                                                                                                                                                                                                                                                            4           ;   /       V        ^�     �   :   <          /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   9   ;          )   signal s1_axis_tlast:  STD_LOGIC:='0';�   8   :          )   signal s1_axis_tvalid: STD_LOGIC:='1';�   7   9          H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�                 <        ����                                                                                                                                                                                                                                                                                                                            4           ;   /       V        ^�     �   ;   <          P   signal s2_axis_tdata  : STD_LOGIC_VECTOR (7 downto 0) := (others=>'0'); --{{{   -   signal s2_axis_tvalid : STD_LOGIC  := '0';   -   signal s2_axis_tlast  : STD_LOGIC  := '0';   3   signal s2_axis_tready : STD_LOGIC  := '1'; --}}}5�_�                 4        ����                                                                                                                                                                                                                                                                                                                            4           ;   /       V        ^�     �   3   <   �    �   4   5   �    5�_�                 @        ����                                                                                                                                                                                                                                                                                                                            <           C   /       V        ^�     �   B   D          /   signal s2_axis_tready: STD_LOGIC:='0'; --}}}�   A   C          )   signal s2_axis_tlast:  STD_LOGIC:='0';�   @   B          )   signal s2_axis_tvalid: STD_LOGIC:='1';�   ?   A          H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�                 <        ����                                                                                                                                                                                                                                                                                                                            <           C   /       V        ^�     �   >   @          )   signal m2_axis_tready: STD_LOGIC:='1';�   =   ?          )   signal m2_axis_tlast:  STD_LOGIC:='0';�   <   >          )   signal m2_axis_tvalid: STD_LOGIC:='0';�   ;   =          M   signal m2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�                 u       ����                                                                                                                                                                                                                                                                                                                            u          x                 ^     �   t   y   �      )           s_axis_tdata  =>m1_axis_tdata,   *           s_axis_tvalid =>m1_axis_tvalid,   )           s_axis_tlast  =>m1_axis_tlast,   *           s_axis_tready =>m1_axis_tready,5�_�                 u       ����                                                                                                                                                                                                                                                                                                                            u          x                 ^     �   t   y   �      )           s_axis_tdata  =>m2_axis_tdata,   *           s_axis_tvalid =>m2_axis_tvalid,   )           s_axis_tlast  =>m2_axis_tlast,   *           s_axis_tready =>m2_axis_tready,5�_�                 q       ����                                                                                                                                                                                                                                                                                                                            t          q                 ^	   % �   p   u   �      )           m_axis_tdata  =>s2_axis_tdata,   *           m_axis_tvalid =>s2_axis_tvalid,   )           m_axis_tlast  =>s2_axis_tlast,   *           m_axis_tready =>s2_axis_tready,5�_�                 }       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^r   & �   |   �   �      )           m_axis_tdata  =>s2_axis_tdata,   *           m_axis_tvalid =>s2_axis_tvalid,   )           m_axis_tlast  =>s2_axis_tlast,   *           m_axis_tready =>s2_axis_tready,5�_�    $             P       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^�     �   O   Q   �      Q            s1_axis_tvalid<= '1'; --que haga de cuentqa que siempre tiene un dato5�_�    &        $   P       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^M     �   O   Q   �      Q            s1_axis_tvalid<= '0'; --que haga de cuentqa que siempre tiene un dato5�_�  $  '  %      &   }       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^�     �   |   �   �      )           m_axis_tdata  =>s1_axis_tdata,   *           m_axis_tvalid =>s1_axis_tvalid,   )           m_axis_tlast  =>s1_axis_tlast,   *           m_axis_tready =>s1_axis_tready,5�_�  &  (          '   <        ����                                                                                                                                                                                                                                                                                                                            }          �                 ^�     �   ;   D   �    �   <   =   �    5�_�  '  )          (   D        ����                                                                                                                                                                                                                                                                                                                            D          G          V       ^�     �   C   D          M   signal m3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{   )   signal m3_axis_tvalid: STD_LOGIC:='0';   )   signal m3_axis_tlast:  STD_LOGIC:='0';   )   signal m3_axis_tready: STD_LOGIC:='1';5�_�  (  *          )   D        ����                                                                                                                                                                                                                                                                                                                            D          G          V       ^�     �   F   H          /   signal s3_axis_tready: STD_LOGIC:='0'; --}}}�   E   G          )   signal s3_axis_tlast:  STD_LOGIC:='0';�   D   F          )   signal s3_axis_tvalid: STD_LOGIC:='1';�   C   E          H   signal s3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�  )  +          *   G   )    ����                                                                                                                                                                                                                                                                                                                            G          G          V       ^�     �   F   H   �      /   signal so_axis_tready: STD_LOGIC:='0'; --}}}5�_�  *  ,          +   D        ����                                                                                                                                                                                                                                                                                                                            D   (       G   (       V   (    ^�     �   F   H   �      )   signal so_axis_tready: STD_LOGIC:='0';�   C   E   �      H   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�  +  -          ,   D        ����                                                                                                                                                                                                                                                                                                                            D   (       G   (       V   (    ^�     �   C   E   �         �   C   E   �    5�_�  ,  .          -   D       ����                                                                                                                                                                                                                                                                                                                            E   (       H   (       V   (    ^      �   C   D             O5�_�  -  /          .   D       ����                                                                                                                                                                                                                                                                                                                            D   (       G   (       V   (    ^   + �   C   E   �    5�_�  .  0          /   E   H    ����                                                                                                                                                                                                                                                                                                                            E   (       H   (       V   (    ^     �   D   F   �      K   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');{{{5�_�  /  1          0   H   )    ����                                                                                                                                                                                                                                                                                                                            E   (       H   (       V   (    ^
     �   G   I   �      /   signal so_axis_tready: STD_LOGIC:='0'; --}}}5�_�  0  2          1   E   (    ����                                                                                                                                                                                                                                                                                                                            H   (       E   (       V   (    ^     �   G   I   �      )   signal so_axis_tready: STD_LOGIC:='0';�   D   F   �      H   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�  1  3          2   E   H    ����                                                                                                                                                                                                                                                                                                                            H   (       E   (       V   (    ^#     �   D   F   �      K   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');{{{5�_�  2  4          3   E   H    ����                                                                                                                                                                                                                                                                                                                            H   (       E   (       V   (    ^$     �   D   F   �      H   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');5�_�  3  7          4   H   *    ����                                                                                                                                                                                                                                                                                                                            E   H       H   /       V   H    ^'     �   G   I   �      /   signal so_axis_tready: STD_LOGIC:='0'; --}}}5�_�  4  8  6      7   F        ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^:     �   G   I   �      *   signal so_axis_tready: STD_LOGIC:='0'; �   E   G   �      )   signal so_axis_tvalid: STD_LOGIC:='1';5�_�  7  9          8   E   I    ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^F     �   D   F   �      I   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0'); 5�_�  8  ;          9   F   )    ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^M   . �   E   G   �      /   signal so_axis_tvalid: STD_LOGIC:='1'; --{{{5�_�  9  <  :      ;   H   &    ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^�     �   G   I   �      0   signal so_axis_tready: STD_LOGIC:='0';  --}}}5�_�  ;  =          <   H   &    ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^�     �   G   I   �      0   signal so_axis_tready: STD_LOGIC:='2';  --}}}5�_�  <  >          =   F   &    ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^�   / �   E   G   �      )   signal so_axis_tvalid: STD_LOGIC:='1';5�_�  =  ?          >   D        ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^�     �   C   D           5�_�  >  @          ?           ����                                                                                                                                                                                                                                                                                                                                      
   *       V   *    ^�     �   	      �      .   signal state   :axiStates := waitingSvalid;�      	   �      architecture arq of all_tb is5�_�  ?  A          @           ����                                                                                                                                                                                                                                                                                                                                      
   *       V   *    ^�     �                 5�_�  @  B          A   )        ����                                                                                                                                                                                                                                                                                                                            )           *           V        ^�     �   (   )          .   signal clk_tb            : STD_LOGIC:= '0';   .   signal rst_tb            : STD_LOGIC:= '0';5�_�  A  C          B           ����                                                                                                                                                                                                                                                                                                                            )           )           V        ^�   0 �   
      �    �         �    5�_�  B  D          C           ����                                                                                                                                                                                                                                                                                                                            +           +           V        ^�     �         �    �         �    5�_�  C  E          D           ����                                                                                                                                                                                                                                                                                                                                       *   "       V        ^�     �   )   +          "   end component split_1to8; --}}}�                    component split_1to8 is --{{{5�_�  D  F          E   �        ����                                                                                                                                                                                                                                                                                                                                       *   "       V        ^�     �   �   �   �    �   �   �   �    5�_�  E  G          F   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^�   1 �   �   �           split_1to8_inst:split_1to8 --{{{5�_�  F  I          G           ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^�   5 �   �   �           split_1to8_inst:split_1to8 --{{{�                "   end component split_1to8; --}}}�                    component split_1to8 is --{{{5�_�  G  J  H      I   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �    �   :   ;   �    5�_�  I  K          J   :   I    ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  J  L          K   :   ,    ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      I   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); -5�_�  K  M          L   :   .    ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      K   signal m1_axis_tdata:  STD_LOGIC_VECTOR (217 downto 0):=(others=>'0'); -5�_�  L  N          M   :   H    ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      J   signal m1_axis_tdata:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0'); -5�_�  M  O          N   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      H   signal m1_axis_tdata:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  N  P          O   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      G   signal m1_axistdata:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  O  Q          P   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      F   signal m1_axisdata:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  P  R          Q   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      E   signal m1_axisata:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  Q  S          R   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      D   signal m1_axista:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  R  T          S   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   9   ;   �      C   signal m1_axisa:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  S  U          T   :       ����                                                                                                                                                                                                                                                                                                                                                             ^+     �   9   :          B   signal m1_axis:  STD_LOGIC_VECTOR (21 downto 0):=(others=>'0');5�_�  T  V          U   R   9    ����                                                                                                                                                                                                                                                                                                                                                             ^+   6 �   Q   S   �      O   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');  --{{{5�_�  U  X          V   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4          9    ^6P   8 �   �   �   �          port map(     )           m_axis_tdata  =>s3_axis_tdata,   *           m_axis_tvalid =>s3_axis_tvalid,   )           m_axis_tlast  =>s3_axis_tlast,   *           m_axis_tready =>s3_axis_tready,   )           s_axis_tdata  =>m3_axis_tdata,   *           s_axis_tvalid =>m3_axis_tvalid,   )           s_axis_tlast  =>m3_axis_tlast,   *           s_axis_tready =>m3_axis_tready,   -           clk           =>clk_tb           ,   4           rst           =>rst_tb           ); --}}}   $slice_2from8_inst:slice_2from8 --{{{       port map(     )           m_axis_tdata  =>s3_axis_tdata,   *           m_axis_tvalid =>s3_axis_tvalid,   )           m_axis_tlast  =>s3_axis_tlast,   *           m_axis_tready =>s3_axis_tready,   )           s_axis_tdata  =>m3_axis_tdata,   *           s_axis_tvalid =>m3_axis_tvalid,   )           s_axis_tlast  =>m3_axis_tlast,   *           s_axis_tready =>m3_axis_tready,   -           clk           =>clk_tb           ,   4           rst           =>rst_tb           ); --}}}�   �   �   �      $slice_1from8_inst:slice_1from8 --{{{5�_�  V  Y  W      X   j        ����                                                                                                                                                                                                                                                                                                                            j          o          V       ^:%     �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      *           m_axis_tready =>so_axis_tready,�   �   �   �      )           m_axis_tlast  =>so_axis_tlast,�   �   �   �      *           m_axis_tvalid =>so_axis_tvalid,�   �   �   �      )           m_axis_tdata  =>so_axis_tdata,�   �   �   �          port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   ~   �   �      %   end process axi_master_proc; --}}}�   }      �            end if;�   |   ~   �               end if;�   {   }   �                  end case;�   z   |   �                        end if;�   y   {   �                           end if;�   x   z   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   w   y   �      .                        s1_axis_tready <= '1';�   v   x   �      .                        m1_axis_tvalid <= '0';�   u   w   �                           else�   t   v   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   s   u   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   r   t   �      Q                     bitCounter := bitCounter+1;                     --incremento�   q   s   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   p   r   �      $               when waitingMready =>�   o   q   �                        end if;�   n   p   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   m   o   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   l   n   �      I                     data           := to_integer(to_signed(data + 1,8));�   k   m   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   j   l   �      )                     bitCounter     := 0;�   i   k   �      +                     s1_axis_tready <= '0';�   h   j   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   g   i   �      $               when waitingSvalid =>�   f   h   �                  case state is�   e   g   �               else�   d   f   �                  data  := 0;�   c   e   �      ,            m1_axis_tdata<= (others => '0');�   b   d   �      !            m1_axis_tvalid<= '0';�   a   c   �      Q            s1_axis_tvalid<= '1'; --que haga de cuentqa que siempre tiene un dato�   `   b   �      !            s1_axis_tready<= '1';�   _   a   �      +            state         <= waitingSvalid;�   ^   `   �               if rst_tb = '0' then�   ]   _   �      !      if rising_edge(clk_tb) then�   \   ^   �         begin�   [   ]   �      2      variable data :integer range -128 to 127:=0;�   Z   \   �      0      variable bitCounter :integer range 0 to 8;�   Y   [   �      ,   axi_master_proc:process (clk_tb) is --{{{�   X   Z   �          rst_tb   <= '1' after 180 ns;�   W   Y   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   T   V   �      0   signal so_axis_tready: STD_LOGIC:='1';  --}}}�   S   U   �      )   signal so_axis_tlast:  STD_LOGIC:='0';�   R   T   �      )   signal so_axis_tvalid: STD_LOGIC:='0';�   Q   S   �      N   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   P   R   �      /   signal s3_axis_tready: STD_LOGIC:='0'; --}}}�   O   Q   �      )   signal s3_axis_tlast:  STD_LOGIC:='0';�   N   P   �      )   signal s3_axis_tvalid: STD_LOGIC:='1';�   M   O   �      H   signal s3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   L   N   �      )   signal m3_axis_tready: STD_LOGIC:='1';�   K   M   �      )   signal m3_axis_tlast:  STD_LOGIC:='0';�   J   L   �      )   signal m3_axis_tvalid: STD_LOGIC:='0';�   I   K   �      M   signal m3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   H   J   �      /   signal s2_axis_tready: STD_LOGIC:='0'; --}}}�   G   I   �      )   signal s2_axis_tlast:  STD_LOGIC:='0';�   F   H   �      )   signal s2_axis_tvalid: STD_LOGIC:='1';�   E   G   �      H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   D   F   �      )   signal m2_axis_tready: STD_LOGIC:='1';�   C   E   �      )   signal m2_axis_tlast:  STD_LOGIC:='0';�   B   D   �      )   signal m2_axis_tvalid: STD_LOGIC:='0';�   A   C   �      M   signal m2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   @   B   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   ?   A   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   >   @   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   =   ?   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   <   >   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   ;   =   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   :   <   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   9   ;   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   i   k          *                     s1_axis_tready<= '0';�   n   p          �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   m   o          o                     m1_axis_tvalid<= '1';                         --como puedo mandar, le avoso que tengo dato�   l   n          J                     data             :=to_integer(to_signed(data + 1,8));�   k   m          I                     m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   j   l          +                     bitCounter       := 0;5�_�  X  Z          Y   j   &    ����                                                                                                                                                                                                                                                                                                                            j          o          V       ^:(   9 �   i   k   �      +                     s1_axis_tready <= '0';5�_�  Y  [          Z   `        ����                                                                                                                                                                                                                                                                                                                            e          `   &       V   &    ^:G   : �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      *           m_axis_tready =>so_axis_tready,�   �   �   �      )           m_axis_tlast  =>so_axis_tlast,�   �   �   �      *           m_axis_tvalid =>so_axis_tvalid,�   �   �   �      )           m_axis_tdata  =>so_axis_tdata,�   �   �   �          port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   ~   �   �      %   end process axi_master_proc; --}}}�   }      �            end if;�   |   ~   �               end if;�   {   }   �                  end case;�   z   |   �                        end if;�   y   {   �                           end if;�   x   z   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   w   y   �      .                        s1_axis_tready <= '1';�   v   x   �      .                        m1_axis_tvalid <= '0';�   u   w   �                           else�   t   v   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   s   u   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   r   t   �      Q                     bitCounter := bitCounter+1;                     --incremento�   q   s   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   p   r   �      $               when waitingMready =>�   o   q   �                        end if;�   n   p   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   m   o   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   l   n   �      I                     data           := to_integer(to_signed(data + 1,8));�   k   m   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   j   l   �      )                     bitCounter     := 0;�   i   k   �      *                     s1_axis_tready <='0';�   h   j   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   g   i   �      $               when waitingSvalid =>�   f   h   �                  case state is�   e   g   �               else�   d   f   �                   data           := 0;�   c   e   �      .            m1_axis_tdata  <= (others => '0');�   b   d   �      "            m1_axis_tvalid <= '0';�   a   c   �      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   `   b   �      "            s1_axis_tready <= '1';�   _   a   �      ,            state          <= waitingSvalid;�   ^   `   �               if rst_tb = '0' then�   ]   _   �      !      if rising_edge(clk_tb) then�   \   ^   �         begin�   [   ]   �      2      variable data :integer range -128 to 127:=0;�   Z   \   �      0      variable bitCounter :integer range 0 to 8;�   Y   [   �      ,   axi_master_proc:process (clk_tb) is --{{{�   X   Z   �          rst_tb   <= '1' after 180 ns;�   W   Y   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   T   V   �      0   signal so_axis_tready: STD_LOGIC:='1';  --}}}�   S   U   �      )   signal so_axis_tlast:  STD_LOGIC:='0';�   R   T   �      )   signal so_axis_tvalid: STD_LOGIC:='0';�   Q   S   �      N   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   P   R   �      /   signal s3_axis_tready: STD_LOGIC:='0'; --}}}�   O   Q   �      )   signal s3_axis_tlast:  STD_LOGIC:='0';�   N   P   �      )   signal s3_axis_tvalid: STD_LOGIC:='1';�   M   O   �      H   signal s3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   L   N   �      )   signal m3_axis_tready: STD_LOGIC:='1';�   K   M   �      )   signal m3_axis_tlast:  STD_LOGIC:='0';�   J   L   �      )   signal m3_axis_tvalid: STD_LOGIC:='0';�   I   K   �      M   signal m3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   H   J   �      /   signal s2_axis_tready: STD_LOGIC:='0'; --}}}�   G   I   �      )   signal s2_axis_tlast:  STD_LOGIC:='0';�   F   H   �      )   signal s2_axis_tvalid: STD_LOGIC:='1';�   E   G   �      H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   D   F   �      )   signal m2_axis_tready: STD_LOGIC:='1';�   C   E   �      )   signal m2_axis_tlast:  STD_LOGIC:='0';�   B   D   �      )   signal m2_axis_tvalid: STD_LOGIC:='0';�   A   C   �      M   signal m2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   @   B   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   ?   A   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   >   @   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   =   ?   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   <   >   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   ;   =   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   :   <   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   9   ;   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   _   a          +            state         <= waitingSvalid;�   d   f                      data  := 0;�   c   e          ,            m1_axis_tdata<= (others => '0');�   b   d          !            m1_axis_tvalid<= '0';�   a   c          Q            s1_axis_tvalid<= '1'; --que haga de cuentqa que siempre tiene un dato�   `   b          !            s1_axis_tready<= '1';5�_�  Z  \          [   �        ����                                                                                                                                                                                                                                                                                                                            e          `   &       V   &    ^Uc     �   �   �   �    �   �   �   �    5�_�  [  ]          \   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^Uj     �   �   �          mapper_inst:mapper --{{{5�_�  \  ^          ]   +        ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^Uo     �   *   :   �    �   +   ,   �    5�_�  ]  _          ^   :        ����                                                                                                                                                                                                                                                                                                                            :           H          V        ^Ur     �   G   I             end component mapper; --}}}�   9   ;             component mapper is --{{{5�_�  ^  `          _   ;        ����                                                                                                                                                                                                                                                                                                                            :           H          V        ^U~     �   :   >   �    �   ;   <   �    5�_�  _  a          `   �       ����                                                                                                                                                                                                                                                                                                                            :           K          V        ^U�     �   �   �   �    �   �   �   �    5�_�  `  b          a   �   
    ����                                                                                                                                                                                                                                                                                                                            :           K          V        ^U�     �   �   �   �         generic(5�_�  a  c          b   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^U�     �   �   �   �      9             N     : natural := 16; --Ancho de la palabra5�_�  b  d          c   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^U�     �   �   �   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto5�_�  c  e          d   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      /             N     := 16; --Ancho de la palabra   ?             ITER  := 10); -- numero de iteraciones por defecto5�_�  d  f          e   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      .             N     = 16; --Ancho de la palabra5�_�  e  g          f   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      >             ITER  = 10); -- numero de iteraciones por defecto5�_�  f  h          g   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �                   N     = 16; 5�_�  g  i          h   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �          port map(  5�_�  h  k          i   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �          port map( 5�_�  i  l  j      k   \        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   [   d   �    �   \   ]   �    5�_�  k  m          l   d        ����                                                                                                                                                                                                                                                                                                                            d           k   /       V        ^U�     �   j   l          /   signal s3_axis_tready: STD_LOGIC:='0'; --}}}�   i   k          )   signal s3_axis_tlast:  STD_LOGIC:='0';�   h   j          )   signal s3_axis_tvalid: STD_LOGIC:='1';�   g   i          H   signal s3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   f   h          )   signal m3_axis_tready: STD_LOGIC:='1';�   e   g          )   signal m3_axis_tlast:  STD_LOGIC:='0';�   d   f          )   signal m3_axis_tvalid: STD_LOGIC:='0';�   c   e          M   signal m3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  l  n          m   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^U�     �   �   �             generic map(                N     = 16;                ITER  = 10);5�_�  m  o          n   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^U�     �   �   �   �    �   �   �   �    5�_�  n  p          o   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      )           m_axis_tdata  =>so_axis_tdata,   *           m_axis_tvalid =>so_axis_tvalid,   )           m_axis_tlast  =>so_axis_tlast,   *           m_axis_tready =>so_axis_tready,5�_�  o  q          p   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      )           m_axis_tdata  =>s1_axis_tdata,   *           m_axis_tvalid =>s1_axis_tvalid,   )           m_axis_tlast  =>s1_axis_tlast,   *           m_axis_tready =>s1_axis_tready,5�_�  p  r          q   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�   ; �   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,   *           s_axis_tvalid =>m1_axis_tvalid,   )           s_axis_tlast  =>m1_axis_tlast,   *           s_axis_tready =>m1_axis_tready,5�_�  q  s          r   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^V     �   �   �   �                   N     = 16;5�_�  r  t          s   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^V   < �   �   �   �                   N     = 16m5�_�  s  u          t   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^V   = �   �   �   �                   ITER  = 10);5�_�  t  v          u   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^V   > �   �   �   �                   ITER  = 10),5�_�  u  w          v   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Vr     �   �   �   �                   N     = 16,                ITER  = 10);5�_�  v  x          w   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Vt     �   �   �   �                   ITER  =>10);�   �   �   �                   N     =>16,5�_�  w  y          x   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Vw   ? �   �   �   �                   ITER  => 10);5�_�  x  z          y   T       ����                                                                                                                                                                                                                                                                                                                            W          T                 ^Z-     �   T   X   �      )   signal m2_axis_tvalid: STD_LOGIC:='0';   )   signal m2_axis_tlast:  STD_LOGIC:='0';   )   signal m2_axis_tready: STD_LOGIC:='1';�   S   U   �      M   signal m2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  y  {          z   T   
    ����                                                                                                                                                                                                                                                                                                                            T   
       W                 ^Z3     �   S   X   �      N   signal m2_axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{   *   signal m2_axis2_tvalid: STD_LOGIC:='0';   *   signal m2_axis2_tlast:  STD_LOGIC:='0';   *   signal m2_axis2_tready: STD_LOGIC:='1';5�_�  z  |          {   X        ����                                                                                                                                                                                                                                                                                                                            X   
       [   
       V   
    ^Z5     �   W   X          H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');   )   signal s2_axis_tvalid: STD_LOGIC:='1';   )   signal s2_axis_tlast:  STD_LOGIC:='0';   /   signal s2_axis_tready: STD_LOGIC:='0'; --}}}5�_�  {  }          |   W   $    ����                                                                                                                                                                                                                                                                                                                            X   
       X   
       V   
    ^Z?     �   V   X   �      '   signal axis2_tready: STD_LOGIC:='1';5�_�  |  ~          }   X        ����                                                                                                                                                                                                                                                                                                                            X   $       g   $       V   $    ^ZF     �   W   X          M   signal m3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{   )   signal m3_axis_tvalid: STD_LOGIC:='0';   )   signal m3_axis_tlast:  STD_LOGIC:='0';   )   signal m3_axis_tready: STD_LOGIC:='1';   H   signal s3_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');   )   signal s3_axis_tvalid: STD_LOGIC:='1';   )   signal s3_axis_tlast:  STD_LOGIC:='0';   /   signal s3_axis_tready: STD_LOGIC:='0'; --}}}   M   signal m4_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{   )   signal m4_axis_tvalid: STD_LOGIC:='0';   )   signal m4_axis_tlast:  STD_LOGIC:='0';   )   signal m4_axis_tready: STD_LOGIC:='1';   H   signal s4_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');   )   signal s4_axis_tvalid: STD_LOGIC:='1';   )   signal s4_axis_tlast:  STD_LOGIC:='0';   /   signal s4_axis_tready: STD_LOGIC:='0'; --}}}5�_�  }            ~   X   
    ����                                                                                                                                                                                                                                                                                                                            X   
       [                 ^ZT     �   W   \   �      N   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{   )   signal so_axis_tvalid: STD_LOGIC:='0';   )   signal so_axis_tlast:  STD_LOGIC:='0';   0   signal so_axis_tready: STD_LOGIC:='1';  --}}}5�_�  ~  �             X       ����                                                                                                                                                                                                                                                                                                                            X          [                 ^ZW     �   X   \   �      &   signal axis_tvalid: STD_LOGIC:='0';   &   signal axis_tlast:  STD_LOGIC:='0';   -   signal axis_tready: STD_LOGIC:='1';  --}}}�   W   Y   �      K   signal axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{5�_�    �          �   X       ����                                                                                                                                                                                                                                                                                                                            X          [                 ^Z\     �   W   \   �      L   signal axiso_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{   '   signal axiso_tvalid: STD_LOGIC:='0';   '   signal axiso_tlast:  STD_LOGIC:='0';   .   signal axiso_tready: STD_LOGIC:='1';  --}}}5�_�  �  �          �   T   E    ����                                                                                                                                                                                                                                                                                                                            X          [                 ^Zc     �   S   U   �      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  �  �          �   T        ����                                                                                                                                                                                                                                                                                                                            T   D       W   '       V   D    ^Zi     �   V   X   �      '   signal axis2_tready: STD_LOGIC:='0';�   S   U   �      E   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');5�_�  �  �          �   T        ����                                                                                                                                                                                                                                                                                                                            T   D       W   '       V   D    ^Zk     �   S   X   �    �   T   U   �    5�_�  �  �          �   X        ����                                                                                                                                                                                                                                                                                                                            X   D       [   '       V   D    ^Zl     �   W   \   �    �   X   Y   �    5�_�  �  �          �   X        ����                                                                                                                                                                                                                                                                                                                            X           [   -       V        ^Zs     �   Z   \          -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   Y   [          '   signal axis2_tlast:  STD_LOGIC:='0';�   X   Z          '   signal axis2_tvalid: STD_LOGIC:='0';�   W   Y          H   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�  �  �          �   \        ����                                                                                                                                                                                                                                                                                                                            \           _   -       V        ^Zz     �   ^   `          -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   ]   _          '   signal axis2_tlast:  STD_LOGIC:='0';�   \   ^          '   signal axis2_tvalid: STD_LOGIC:='0';�   [   ]          H   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   �   �   �      )           m_axis_tdata  =>s2_axis_tdata,   *           m_axis_tvalid =>s2_axis_tvalid,   )           m_axis_tlast  =>s2_axis_tlast,   *           m_axis_tready =>s2_axis_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   �   �   �      '           m_axis_tvalid =>axis_tvalid,   &           m_axis_tlast  =>axis_tlast,   '           m_axis_tready =>axis_tready,�   �   �   �      &           m_axis_tdata  =>axis_tdata,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   �   �   �      )           s_axis_tdata  =>m2_axis_tdata,   *           s_axis_tvalid =>m2_axis_tvalid,   )           s_axis_tlast  =>m2_axis_tlast,   *           s_axis_tready =>m2_axis_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   �   �   �      '           s_axis_tvalid =>axis_tvalid,   &           s_axis_tlast  =>axis_tlast,   '           s_axis_tready =>axis_tready,�   �   �   �      &           s_axis_tdata  =>axis_tdata,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   �   �   �      )           m_axis_tdata  =>so_axis_tdata,   *           m_axis_tvalid =>so_axis_tvalid,   )           m_axis_tlast  =>so_axis_tlast,   *           m_axis_tready =>so_axis_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�   @ �   �   �   �      '           m_axis_tvalid =>axis_tvalid,   &           m_axis_tlast  =>axis_tlast,   '           m_axis_tready =>axis_tready,�   �   �   �      &           m_axis_tdata  =>axis_tdata,5�_�  �  �          �   T   E    ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   S   U   �      H   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�  �  �          �   X   E    ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   W   Y   �      H   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�  �  �          �   X   E    ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   W   Y   �      J   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');--{{{5�_�  �  �          �   \   E    ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   [   ]   �      H   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');{{{5�_�  �  �          �   c   G    ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�     �   c   e   �    5�_�  �  �          �   e        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^Z�   B �   d   e           5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^��   C �   �   �   �                   ITER  => 10)5�_�  �  �          �   z   0    ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�E     �   z   |   �                           �   z   |   �    5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�M     �   z   |   �                           if(5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�O     �   z   |   �                           if(5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�O     �   z   }   �                           if5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�Z     �   {   |           5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�[     �   {   }   �    �   |   }   �    5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�]     �   |      �                           �   |   ~   �    5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�f     �   |   ~   �                        else if5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�f     �   |   ~   �                        ele if5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�f     �   |   ~   �                        el if5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�h     �   |   ~   �                        elif5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�m     �   |   ~   �                           else if5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�n     �   }      �                              �   }      �    5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�t     �   }      �    �   ~      �    5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�u     �   }      �      %                     if data<127 then5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�}     �   }      �      (                        if data<127 then5�_�  �  �          �   ~   "    ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^�~     �   }      �      (                        if data>127 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^��     �   z   |   �      %                     if data<127 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^��     �   z   |   �      %                     if data-127 then5�_�  �  �          �   {        ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^��     �   z   {          %                     if data=127 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^��     �   z   |   �    �   {   |   �    5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^��     �   {   }   �    �   |   }   �    5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^��     �   {   }   �      I                     data           := to_integer(to_signed(data + 1,8));5�_�  �  �          �   |   *    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^��     �   {   }   �      L                        data           := to_integer(to_signed(data + 1,8));5�_�  �  �          �   |   .    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^��     �   {   }   �      P                        data           := -128to_integer(to_signed(data + 1,8));5�_�  �  �          �   |   .    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^��     �   |   ~   �                              �   |   ~   �    5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            ~          ~          V       ^��     �   }             I                     data           := to_integer(to_signed(data + 1,8));5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                      �          V       ^��     �   ~                                  else   (                        if data>128 then                           5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                V       ^��     �   ~              5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^��     �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      (           s_axis_tready =>axis2_tready,�   �   �   �      '           s_axis_tlast  =>axis2_tlast,�   �   �   �      (           s_axis_tvalid =>axis2_tvalid,�   �   �   �      '           s_axis_tdata  =>axis2_tdata,�   �   �   �      (           m_axis_tready =>axisO_tready,�   �   �   �      '           m_axis_tlast  =>axisO_tlast,�   �   �   �      (           m_axis_tvalid =>axisO_tvalid,�   �   �   �      '           m_axis_tdata  =>axisO_tdata,�   �   �   �          port map(  �   �   �   �                   ITER  => 5)�   �   �   �                   N     => 16,�   �   �   �         generic map(�   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      (           m_axis_tready =>axis2_tready,�   �   �   �      '           m_axis_tlast  =>axis2_tlast,�   �   �   �      (           m_axis_tvalid =>axis2_tvalid,�   �   �   �      '           m_axis_tdata  =>axis2_tdata,�   �   �   �          port map(�   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      %   end process axi_master_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end if;�   �   �   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                        s1_axis_tready <= '1';�   �   �   �      .                        m1_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   �   �   �      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   �   �   �                        end if;�   �   �   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�      �   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   ~   �   �      I                     data           := to_integer(to_signed(data + 1,8));�   }      �      L                        data           := to_integer(to_signed(data + 1,8));�   |   ~   �                           else�   {   }   �      /                        data           := -128;�   z   |   �      %                     if data=127 then�   y   {   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   x   z   �      )                     bitCounter     := 0;�   w   y   �      *                     s1_axis_tready <='0';�   v   x   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingSvalid =>�   t   v   �                  case state is�   s   u   �               else�   r   t   �                   data           := 0;�   q   s   �      .            m1_axis_tdata  <= (others => '0');�   p   r   �      "            m1_axis_tvalid <= '0';�   o   q   �      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   n   p   �      "            s1_axis_tready <= '1';�   m   o   �      ,            state          <= waitingSvalid;�   l   n   �               if rst_tb = '0' then�   k   m   �      !      if rising_edge(clk_tb) then�   j   l   �         begin�   i   k   �      2      variable data :integer range -128 to 127:=0;�   h   j   �      0      variable bitCounter :integer range 0 to 8;�   g   i   �      ,   axi_master_proc:process (clk_tb) is --{{{�   f   h   �          rst_tb   <= '1' after 180 ns;�   e   g   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   b   d   �      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   a   c   �      '   signal axisO_tlast:  STD_LOGIC:='0';�   `   b   �      '   signal axisO_tvalid: STD_LOGIC:='0';�   _   a   �      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   ^   `   �      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   ]   _   �      '   signal axis4_tlast:  STD_LOGIC:='0';�   \   ^   �      '   signal axis4_tvalid: STD_LOGIC:='0';�   [   ]   �      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   Z   \   �      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   Y   [   �      '   signal axis3_tlast:  STD_LOGIC:='0';�   X   Z   �      '   signal axis3_tvalid: STD_LOGIC:='0';�   W   Y   �      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   V   X   �      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   U   W   �      '   signal axis2_tlast:  STD_LOGIC:='0';�   T   V   �      '   signal axis2_tvalid: STD_LOGIC:='0';�   S   U   �      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   R   T   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   Q   S   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   P   R   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   O   Q   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   N   P   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   M   O   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   L   N   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   K   M   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   J   L   �         end component cordic; --}}}�   I   K   �      *           rst           : in  STD_LOGIC);�   H   J   �      )           clk           : in  STD_LOGIC;�   F   H   �      )           s_axis_tready : out STD_LOGIC;�   E   G   �      )           s_axis_tlast  : in  STD_LOGIC;�   D   F   �      )           s_axis_tvalid : in  STD_LOGIC;�   C   E   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C   �      )           m_axis_tready : in  STD_LOGIC;�   @   B   �      )           m_axis_tlast  : out STD_LOGIC;�   ?   A   �      )           m_axis_tvalid : out STD_LOGIC;�   >   @   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?   �      	    port(�   <   >   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =   �      9             N     : natural := 16; --Ancho de la palabra�   :   <   �         generic(�   9   ;   �         component cordic is --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   {   }          /                        data           := -128;5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            |           |           V        ^��     �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      (           s_axis_tready =>axis2_tready,�   �   �   �      '           s_axis_tlast  =>axis2_tlast,�   �   �   �      (           s_axis_tvalid =>axis2_tvalid,�   �   �   �      '           s_axis_tdata  =>axis2_tdata,�   �   �   �      (           m_axis_tready =>axisO_tready,�   �   �   �      '           m_axis_tlast  =>axisO_tlast,�   �   �   �      (           m_axis_tvalid =>axisO_tvalid,�   �   �   �      '           m_axis_tdata  =>axisO_tdata,�   �   �   �          port map(  �   �   �   �                   ITER  => 5)�   �   �   �                   N     => 16,�   �   �   �         generic map(�   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      (           m_axis_tready =>axis2_tready,�   �   �   �      '           m_axis_tlast  =>axis2_tlast,�   �   �   �      (           m_axis_tvalid =>axis2_tvalid,�   �   �   �      '           m_axis_tdata  =>axis2_tdata,�   �   �   �          port map(�   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      %   end process axi_master_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end if;�   �   �   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                        s1_axis_tready <= '1';�   �   �   �      .                        m1_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   �   �   �      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   �   �   �                        end if;�   �   �   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�      �   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   ~   �   �      I                     data           := to_integer(to_signed(data + 1,8));�   }      �      L                        data           := to_integer(to_signed(data + 1,8));�   |   ~   �                           else�   {   }   �      /                        data           := -128;�   z   |   �      %                     if data=127 then�   y   {   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   x   z   �      )                     bitCounter     := 0;�   w   y   �      *                     s1_axis_tready <='0';�   v   x   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingSvalid =>�   t   v   �                  case state is�   s   u   �               else�   r   t   �                   data           := 0;�   q   s   �      .            m1_axis_tdata  <= (others => '0');�   p   r   �      "            m1_axis_tvalid <= '0';�   o   q   �      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   n   p   �      "            s1_axis_tready <= '1';�   m   o   �      ,            state          <= waitingSvalid;�   l   n   �               if rst_tb = '0' then�   k   m   �      !      if rising_edge(clk_tb) then�   j   l   �         begin�   i   k   �      2      variable data :integer range -128 to 127:=0;�   h   j   �      0      variable bitCounter :integer range 0 to 8;�   g   i   �      ,   axi_master_proc:process (clk_tb) is --{{{�   f   h   �          rst_tb   <= '1' after 180 ns;�   e   g   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   b   d   �      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   a   c   �      '   signal axisO_tlast:  STD_LOGIC:='0';�   `   b   �      '   signal axisO_tvalid: STD_LOGIC:='0';�   _   a   �      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   ^   `   �      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   ]   _   �      '   signal axis4_tlast:  STD_LOGIC:='0';�   \   ^   �      '   signal axis4_tvalid: STD_LOGIC:='0';�   [   ]   �      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   Z   \   �      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   Y   [   �      '   signal axis3_tlast:  STD_LOGIC:='0';�   X   Z   �      '   signal axis3_tvalid: STD_LOGIC:='0';�   W   Y   �      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   V   X   �      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   U   W   �      '   signal axis2_tlast:  STD_LOGIC:='0';�   T   V   �      '   signal axis2_tvalid: STD_LOGIC:='0';�   S   U   �      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   R   T   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   Q   S   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   P   R   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   O   Q   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   N   P   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   M   O   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   L   N   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   K   M   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   J   L   �         end component cordic; --}}}�   I   K   �      *           rst           : in  STD_LOGIC);�   H   J   �      )           clk           : in  STD_LOGIC;�   F   H   �      )           s_axis_tready : out STD_LOGIC;�   E   G   �      )           s_axis_tlast  : in  STD_LOGIC;�   D   F   �      )           s_axis_tvalid : in  STD_LOGIC;�   C   E   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C   �      )           m_axis_tready : in  STD_LOGIC;�   @   B   �      )           m_axis_tlast  : out STD_LOGIC;�   ?   A   �      )           m_axis_tvalid : out STD_LOGIC;�   >   @   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?   �      	    port(�   <   >   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =   �      9             N     : natural := 16; --Ancho de la palabra�   :   <   �         generic(�   9   ;   �         component cordic is --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   {   }          /                        data           := -128;5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            |           |           V        ^��     �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      (           s_axis_tready =>axis2_tready,�   �   �   �      '           s_axis_tlast  =>axis2_tlast,�   �   �   �      (           s_axis_tvalid =>axis2_tvalid,�   �   �   �      '           s_axis_tdata  =>axis2_tdata,�   �   �   �      (           m_axis_tready =>axisO_tready,�   �   �   �      '           m_axis_tlast  =>axisO_tlast,�   �   �   �      (           m_axis_tvalid =>axisO_tvalid,�   �   �   �      '           m_axis_tdata  =>axisO_tdata,�   �   �   �          port map(  �   �   �   �                   ITER  => 5)�   �   �   �                   N     => 16,�   �   �   �         generic map(�   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      (           m_axis_tready =>axis2_tready,�   �   �   �      '           m_axis_tlast  =>axis2_tlast,�   �   �   �      (           m_axis_tvalid =>axis2_tvalid,�   �   �   �      '           m_axis_tdata  =>axis2_tdata,�   �   �   �          port map(�   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      %   end process axi_master_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end if;�   �   �   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                        s1_axis_tready <= '1';�   �   �   �      .                        m1_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   �   �   �      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   �   �   �                        end if;�   �   �   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�      �   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   ~   �   �      I                     data           := to_integer(to_signed(data + 1,8));�   }      �      L                        data           := to_integer(to_signed(data + 1,8));�   |   ~   �                           else�   {   }   �      %                        data := -128;�   z   |   �      %                     if data=127 then�   y   {   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   x   z   �      )                     bitCounter     := 0;�   w   y   �      *                     s1_axis_tready <='0';�   v   x   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingSvalid =>�   t   v   �                  case state is�   s   u   �               else�   r   t   �                   data           := 0;�   q   s   �      .            m1_axis_tdata  <= (others => '0');�   p   r   �      "            m1_axis_tvalid <= '0';�   o   q   �      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   n   p   �      "            s1_axis_tready <= '1';�   m   o   �      ,            state          <= waitingSvalid;�   l   n   �               if rst_tb = '0' then�   k   m   �      !      if rising_edge(clk_tb) then�   j   l   �         begin�   i   k   �      2      variable data :integer range -128 to 127:=0;�   h   j   �      0      variable bitCounter :integer range 0 to 8;�   g   i   �      ,   axi_master_proc:process (clk_tb) is --{{{�   f   h   �          rst_tb   <= '1' after 180 ns;�   e   g   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   b   d   �      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   a   c   �      '   signal axisO_tlast:  STD_LOGIC:='0';�   `   b   �      '   signal axisO_tvalid: STD_LOGIC:='0';�   _   a   �      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   ^   `   �      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   ]   _   �      '   signal axis4_tlast:  STD_LOGIC:='0';�   \   ^   �      '   signal axis4_tvalid: STD_LOGIC:='0';�   [   ]   �      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   Z   \   �      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   Y   [   �      '   signal axis3_tlast:  STD_LOGIC:='0';�   X   Z   �      '   signal axis3_tvalid: STD_LOGIC:='0';�   W   Y   �      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   V   X   �      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   U   W   �      '   signal axis2_tlast:  STD_LOGIC:='0';�   T   V   �      '   signal axis2_tvalid: STD_LOGIC:='0';�   S   U   �      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   R   T   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   Q   S   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   P   R   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   O   Q   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   N   P   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   M   O   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   L   N   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   K   M   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   J   L   �         end component cordic; --}}}�   I   K   �      *           rst           : in  STD_LOGIC);�   H   J   �      )           clk           : in  STD_LOGIC;�   F   H   �      )           s_axis_tready : out STD_LOGIC;�   E   G   �      )           s_axis_tlast  : in  STD_LOGIC;�   D   F   �      )           s_axis_tvalid : in  STD_LOGIC;�   C   E   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C   �      )           m_axis_tready : in  STD_LOGIC;�   @   B   �      )           m_axis_tlast  : out STD_LOGIC;�   ?   A   �      )           m_axis_tvalid : out STD_LOGIC;�   >   @   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?   �      	    port(�   <   >   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =   �      9             N     : natural := 16; --Ancho de la palabra�   :   <   �         generic(�   9   ;   �         component cordic is --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   {   }          /                        data           := -128;5�_�  �  �          �   ~        ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^��   D �   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      (           s_axis_tready =>axis2_tready,�   �   �   �      '           s_axis_tlast  =>axis2_tlast,�   �   �   �      (           s_axis_tvalid =>axis2_tvalid,�   �   �   �      '           s_axis_tdata  =>axis2_tdata,�   �   �   �      (           m_axis_tready =>axisO_tready,�   �   �   �      '           m_axis_tlast  =>axisO_tlast,�   �   �   �      (           m_axis_tvalid =>axisO_tvalid,�   �   �   �      '           m_axis_tdata  =>axisO_tdata,�   �   �   �          port map(  �   �   �   �                   ITER  => 5)�   �   �   �                   N     => 16,�   �   �   �         generic map(�   �   �   �      4           rst           =>rst_tb           ); --}}}�   �   �   �      -           clk           =>clk_tb           ,�   �   �   �      *           s_axis_tready =>m1_axis_tready,�   �   �   �      )           s_axis_tlast  =>m1_axis_tlast,�   �   �   �      *           s_axis_tvalid =>m1_axis_tvalid,�   �   �   �      )           s_axis_tdata  =>m1_axis_tdata,�   �   �   �      (           m_axis_tready =>axis2_tready,�   �   �   �      '           m_axis_tlast  =>axis2_tlast,�   �   �   �      (           m_axis_tvalid =>axis2_tvalid,�   �   �   �      '           m_axis_tdata  =>axis2_tdata,�   �   �   �          port map(�   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      6--           rst           =>rst_tb           ); --}}}�   �   �   �      /--           clk           =>clk_tb           ,�   �   �   �      ,--           s_axis_tready =>m3_axis_tready,�   �   �   �      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �   �      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �   �      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �   �      ,--           m_axis_tready =>s3_axis_tready,�   �   �   �      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �   �      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �   �      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �   �      --    port map(  �   �   �   �      %   end process axi_master_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end if;�   �   �   �      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                        s1_axis_tready <= '1';�   �   �   �      .                        m1_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   �   �   �      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �   �      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   �   �   �                        end if;�   �   �   �      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�      �   �      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   ~   �   �      I                     data           := to_integer(to_signed(data + 1,8));�   }      �      B                        data := to_integer(to_signed(data + 1,8));�   |   ~   �                           else�   {   }   �      %                        data := -128;�   z   |   �      %                     if data=127 then�   y   {   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   x   z   �      )                     bitCounter     := 0;�   w   y   �      *                     s1_axis_tready <='0';�   v   x   �      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingSvalid =>�   t   v   �                  case state is�   s   u   �               else�   r   t   �                   data           := 0;�   q   s   �      .            m1_axis_tdata  <= (others => '0');�   p   r   �      "            m1_axis_tvalid <= '0';�   o   q   �      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   n   p   �      "            s1_axis_tready <= '1';�   m   o   �      ,            state          <= waitingSvalid;�   l   n   �               if rst_tb = '0' then�   k   m   �      !      if rising_edge(clk_tb) then�   j   l   �         begin�   i   k   �      2      variable data :integer range -128 to 127:=0;�   h   j   �      0      variable bitCounter :integer range 0 to 8;�   g   i   �      ,   axi_master_proc:process (clk_tb) is --{{{�   f   h   �          rst_tb   <= '1' after 180 ns;�   e   g   �      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   b   d   �      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   a   c   �      '   signal axisO_tlast:  STD_LOGIC:='0';�   `   b   �      '   signal axisO_tvalid: STD_LOGIC:='0';�   _   a   �      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   ^   `   �      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   ]   _   �      '   signal axis4_tlast:  STD_LOGIC:='0';�   \   ^   �      '   signal axis4_tvalid: STD_LOGIC:='0';�   [   ]   �      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   Z   \   �      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   Y   [   �      '   signal axis3_tlast:  STD_LOGIC:='0';�   X   Z   �      '   signal axis3_tvalid: STD_LOGIC:='0';�   W   Y   �      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   V   X   �      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   U   W   �      '   signal axis2_tlast:  STD_LOGIC:='0';�   T   V   �      '   signal axis2_tvalid: STD_LOGIC:='0';�   S   U   �      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   R   T   �      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   Q   S   �      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   P   R   �      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   O   Q   �      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   N   P   �      )   signal m1_axis_tready: STD_LOGIC:='1';�   M   O   �      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   L   N   �      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   K   M   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   J   L   �         end component cordic; --}}}�   I   K   �      *           rst           : in  STD_LOGIC);�   H   J   �      )           clk           : in  STD_LOGIC;�   F   H   �      )           s_axis_tready : out STD_LOGIC;�   E   G   �      )           s_axis_tlast  : in  STD_LOGIC;�   D   F   �      )           s_axis_tvalid : in  STD_LOGIC;�   C   E   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C   �      )           m_axis_tready : in  STD_LOGIC;�   @   B   �      )           m_axis_tlast  : out STD_LOGIC;�   ?   A   �      )           m_axis_tvalid : out STD_LOGIC;�   >   @   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?   �      	    port(�   <   >   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =   �      9             N     : natural := 16; --Ancho de la palabra�   :   <   �         generic(�   9   ;   �         component cordic is --{{{�   8   :   �         end component mapper; --}}}�   7   9   �      *           rst           : in  STD_LOGIC);�   6   8   �      )           clk           : in  STD_LOGIC;�   4   6   �      )           s_axis_tready : out STD_LOGIC;�   3   5   �      )           s_axis_tlast  : in  STD_LOGIC;�   2   4   �      )           s_axis_tvalid : in  STD_LOGIC;�   1   3   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1   �      )           m_axis_tready : in  STD_LOGIC;�   .   0   �      )           m_axis_tlast  : out STD_LOGIC;�   -   /   �      )           m_axis_tvalid : out STD_LOGIC;�   ,   .   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -   �      	    port(�   *   ,   �         component mapper is --{{{�   )   +   �      $   end component slice_2from8; --}}}�   (   *   �      *           rst           : in  STD_LOGIC);�   '   )   �      )           clk           : in  STD_LOGIC;�   %   '   �      )           s_axis_tready : out STD_LOGIC;�   $   &   �      )           s_axis_tlast  : in  STD_LOGIC;�   #   %   �      )           s_axis_tvalid : in  STD_LOGIC;�   "   $   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "   �      )           m_axis_tready : in  STD_LOGIC;�      !   �      )           m_axis_tlast  : out STD_LOGIC;�          �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_2from8 is --{{{�         �      $   end component slice_1from8; --}}}�         �      *           rst           : in  STD_LOGIC);�         �      )           clk           : in  STD_LOGIC;�         �      )           s_axis_tready : out STD_LOGIC;�         �      )           s_axis_tlast  : in  STD_LOGIC;�         �      )           s_axis_tvalid : in  STD_LOGIC;�         �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      )           m_axis_tready : in  STD_LOGIC;�         �      )           m_axis_tlast  : out STD_LOGIC;�         �      )           m_axis_tvalid : out STD_LOGIC;�         �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         �      	    port(�         �      "   component slice_1from8 is --{{{�         �      .   signal rst_tb            : STD_LOGIC:= '0';�   
      �      .   signal clk_tb            : STD_LOGIC:= '0';�      
   �      4   signal state   :axiStates := waitingSvalid; --}}}�      	   �      6   type   axiStates is (waitingSvalid, waitingMready);�   }             L                        data           := to_integer(to_signed(data + 1,8));5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^�   E �   ~             I                     data           := to_integer(to_signed(data + 1,8));5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^�   G �   ~   �   �                              �   ~   �   �    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^�   H �   ~   �   �                           end if5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^��   I �   z   |   �      %                     if data=127 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^�7     �   z   |   �      %                     if data=120 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            ~           ~           V        ^�8   K �   z   |   �      %                     if data=128 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            {                           ^��     �   {   �   �      %                        data := -128;                        else   B                        data := to_integer(to_signed(data + 1,8));                        end if;�   z   |   �      %                     if data=127 then5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            {                           ^��     �   z   |   �    �   {   |   �    5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      '                     --   data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      &                     -   data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      %                        data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      $                       data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      #                      data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      "                     data := -128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      #                     data := 1-128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      "                     data := 1128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��     �   z   |   �      !                     data := 128;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��   M �   z   |   �                            data := 18;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^��   N �   z   |   �                           data := 1;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^�-     �   z   |   �                           data := 0;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^�.   O �   z   |   �      !                     data := 140;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^     �   �   �   �                   ITER  => 5)5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^   P �   �   �   �                   ITER  => 105)5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^+   Q �   z   |   �                            data := 14;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^k   R �   z   |   �                           data := 1;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^     �   z   |   �                           data := 0;5�_�  �  �          �   {       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^   S �   z   |   �                           data := 1;5�_�  �  �          �   j       ����                                                                                                                                                                                                                                                                                                                            |          �                 ^Q     �   i   k   �    �   j   k   �    5�_�  �  �          �   j       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^S     �   i   k   �      2      variable data :integer range -128 to 127:=0;5�_�  �  �          �   k       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^U     �   j   l   �      2      variable data :integer range -128 to 127:=0;5�_�  �  �          �   t       ����                                                                                                                                                                                                                                                                                                                            }          �                 ^Z     �   s   u   �    �   t   u   �    5�_�  �  �          �   t       ����                                                                                                                                                                                                                                                                                                                            ~          �                 ^[     �   s   u   �                   data           := 0;5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                            ~          �                 ^]     �   t   v   �                   data           := 0;5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                            ~          �                 ^_     �   t   v   �                   data2          := 0;5�_�  �  �          �   t       ����                                                                                                                                                                                                                                                                                                                            ~          �                 ^`     �   s   u   �      !            data1           := 0;5�_�  �  �          �   t       ����                                                                                                                                                                                                                                                                                                                            ~          �                 ^a     �   s   u   �                   data1          := 0;5�_�  �  �          �   }        ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^h     �   |   }                               data := 3;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^h     �   {   }   �    �   |   }   �    5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            ~          ~          V       ^i     �   {   }   �                           data := 3;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            ~          ~          V       ^m     �   {   }   �                            data1 := 3;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            ~          ~          V       ^n     �   {   }   �      !                     data1 := 13;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            ~          ~          V       ^q     �   {   }   �    �   |   }   �    5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                                                V       ^r     �   {   }   �                            data1 := 1;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                                                V       ^t     �   {   }   �                            data2 := 1;5�_�  �  �          �   |        ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^u     �   {   |                                data2 := 0;5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^v     �   |   ~   �    �   }   ~   �    5�_�  �  �          �   ~   F    ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^x     �   }      �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^|   U �   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^�     �   {   }   �                            data1 := 1;5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^�   V �   |   ~   �                            data2 := 0;5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^     �   �   �   �      M                        m1_axis_tdata<= std_logic_vector(to_signed(data2,8));5�_�  �  �          �   ~   F    ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^     �   }      �      L                     m1_axis_tdata  <= std_logic_vector(to_signed(data1,8));5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^!     �   {   }   �                            data1 := 0;5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^"     �   |   }                                data2 := 1;5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^$     �   t   v   �                  data2         := 0;5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                            |          |          V       ^'     �   t   u          "            data2    sfdd    := 0;5�_�  �  �          �   t       ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^(     �   s   u   �                  data1         := 0;5�_�  �  �          �   j       ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^+     �   i   k   �      3      variable data1 :integer range -128 to 127:=0;5�_�  �  �          �   k       ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^,   W �   j   k          2      variable data2:integer range -128 to 127:=0;5�_�  �  �          �   �   G    ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^B   X �   �   �   �      M                        m1_axis_tdata<= std_logic_vector(to_signed(data1,8));5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^M     �   {   }   �      '                     --if data=127 then5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^N     �   {   }   �      &                     -if data=127 then5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^O     �   {   }   �      %                     if data=127 then5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^Y     �   |   ~   �      '                     --   data := -128;5�_�  �  �          �   }       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^Y     �   |   ~   �      &                     -   data := -128;5�_�  �  �          �   z       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^_     �   y   {   �                           data := 0;5�_�  �  �          �   |       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^c     �   {   }   �      #                     if data=0 then5�_�  �  �          �   }        ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^e     �   |   ~   �      %                        data := -128;5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^g     �   }      �                           --else5�_�  �  �          �   ~       ����                                                                                                                                                                                                                                                                                                                            z          z          V       ^g     �   }      �                           -else5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                V       ^k     �   ~   �   �    �      �   �    �   ~             D                     --   data := to_integer(to_signed(data + 1,8));5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                          !       V       ^m     �   ~   �   �      "                        data := 0;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                          !       V       ^o     �      �   �                           --end if;5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                          !       V       ^o   Y �      �   �                           -end if;5�_�  �             �   z       ����                                                                                                                                                                                                                                                                                                                                          !       V       ^�     �   y   z                               data := 1;5�_�  �                s       ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�   [ �   r   t   �                  data         := 0;5�_�                  j   0    ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^f     �   i   k   �      2      variable data :integer range -128 to 127:=0;5�_�                 s        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^k   \ �   r   t   �                  data         := 1;5�_�                 ~        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^{   ] �   }      �      "                        data := 1;5�_�                 {       ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^     �   z   |   �      #                     if data=1 then5�_�                 |        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   {   }   �      "                        data := 0;5�_�                 ~        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�   ^ �   }      �      "                        data := 2;5�_�                 {       ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   z   |   �      #                     if data=0 then5�_�    	             s        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   r   t   �       --            data         := 1;5�_�    
          	   s        ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   r   t   �      -            data         := 1;5�_�  	            
   j   0    ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   i   k   �      2      variable data :integer range -128 to 127:=1;5�_�  
               {       ����                                                                                                                                                                                                                                                                                                                            ~           ~   !       V       ^�     �   z   |   �      #                     if data=2 then5�_�                 {        ����                                                                                                                                                                                                                                                                                                                            {          ~          V       ^�     �   z   {          #                     if data=0 then   "                        data := 2;                        else   "                        data := 0;5�_�                 z       ����                                                                                                                                                                                                                                                                                                                            {          {          V       ^�     �   y   ~   �    �   z   {   �    5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �   ~                                  end if;5�_�                 ~       ����                                                                                                                                                                                                                                                                                                                                                V       ^�     �   }      �    �   ~      �    5�_�                 s       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^�   _ �   r   t   �                  data         := 1;5�_�                 {        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^�   ` �   z   |   �      "                        data := 2;5�_�               j   1    ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^     �   i   k   �    �   j   k   �    5�_�                 k       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^     �   j   l   �      2      variable data :integer range -128 to 127:=0;5�_�                 k       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^      �   j   l   �      3      variable data1 :integer range -128 to 127:=0;5�_�                 k   '    ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^'     �   j   l   �      <      variable data1 :std_logic_vector range -128 to 127:=0;5�_�                 k   3    ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^-     �   j   l   �      H      variable data1 :std_logic_vector (3 downto 0)range -128 to 127:=0;5�_�                 {       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^5     �   z   |   �      #                     if data=0 then5�_�                 {       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^7     �   z   |   �      %                     if data=150 then5�_�                 |        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^8     �   {   }   �      "                        data := 3;5�_�                 }        ����                                                                                                                                                                                                                                                                                                                            }          ~           V        ^:     �   |   }                               else   "                        data := 0;5�_�                 ~   .    ����                                                                                                                                                                                                                                                                                                                            }          }           V        ^=     �   }      �    �   ~      �    5�_�                 ~       ����                                                                                                                                                                                                                                                                                                                            }          }           V        ^>     �   }      �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                    '    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^E     �   ~   �   �      K                     m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                     +    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^F     �   ~   �   �      0                     m1_axis_tdata  <= data,8));5�_�    !                 8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^L     �   ~   �   �      =                     m1_axis_tdata  <= data1(1 downto 0),8));5�_�     "          !      8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^L     �   ~   �   �      <                     m1_axis_tdata  <= data1(1 downto 0)8));5�_�  !  #          "      8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^M     �   ~   �   �      ;                     m1_axis_tdata  <= data1(1 downto 0)));5�_�  "  $          #      8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^N     �   ~   �   �      :                     m1_axis_tdata  <= data1(1 downto 0));5�_�  #  %          $   �   %    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^T     �   �   �   �      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   5�_�  $  &          %   �   0    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^X     �   �   �   �    �   �   �   �    5�_�  %  '          &   �       ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^[     �   �   �   �      L                        m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�  &  (          '   �       ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^\     �   �   �   �      9                     m1_axis_tdata  <= data1(1 downto 0);5�_�  '  )          (   �   0    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^^     �   �   �   �      <                        m1_axis_tdata  <= data1(1 downto 0);5�_�  (  *          )   �   9    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^_     �   �   �   �      <                        m1_axis_tdata  <= data1(3 downto 0);5�_�  )  +          *   �   8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^a     �   �   �   �      <                        m1_axis_tdata  <= data1(3 downto 1);5�_�  *  ,          +   �   8    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^c     �   �   �   �      <                        m1_axis_tdata  <= data1(3 downtol1);5�_�  +  -          ,   �   9    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^c     �   �   �   �      <                        m1_axis_tdata  <= data1(3 downto 1);5�_�  ,  .          -   |   !    ����                                                                                                                                                                                                                                                                                                                               '          A       v   A    ^l   a �   |      �                              �   |   ~   �    5�_�  -  /          .   {       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^}     �   z   |   �      $                     if data=15 then5�_�  .  0          /   |       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^~     �   {   }   �      "                        data := 0;5�_�  /  1          0   ~       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   }      �      )                        data := data + 1;5�_�  0  2          1   ~   %    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   }      �      *                        data1 := data + 1;5�_�  1  3          2   {       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   z   |   �      %                     if data1=15 then5�_�  2  4          3   |       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   {   }   �      #                        data1 := 0;5�_�  3  5          4   ~       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   }      �      +                        data1 := data1 + 1;5�_�  4  6          5   ~   %    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   }      �      +                        data2 := data1 + 1;5�_�  5  7          6   k       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   j   l   �    �   k   l   �    5�_�  6  8          7   l       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   k   m   �      4      variable data1 :std_logic_vector (3 downto 0);5�_�  7  9          8   l       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   k   m   �      4      variable data2 :std_logic_vector (3 downto 0);5�_�  8  :          9   l       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   k   m   �      +      variable data2 :natural (3 downto 0);5�_�  9  <          :   l   +    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   k   m   �      8      variable data2 :natural range 0 to 15(3 downto 0);5�_�  :  =  ;      <   �       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   �   �   �                           �   �   �   �    5�_�  <  >          =   �       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   �   �   �      3                     data1 := to_unsigned(data2,4);5�_�  =  ?          >   �   C    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�   b �   �   �   �      D                     data1 := std_logic_vector(to_unsigned(data2,4);5�_�  >  @          ?   �   '    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�   c �   �   �   �      9                     m1_axis_tdata  <= data1(1 downto 0);5�_�  ?  A          @   �   *    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^
   d �   �   �   �      <                        m1_axis_tdata  <= data1(3 downto 2);5�_�  @  H          A   �   '    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^   e �   �   �   �      A                     m1_axis_tdata  <= x"00" & data1(1 downto 0);5�_�  A  I  B      H   �   *    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^@   g �   �   �   �      @                     m1_axis_tdata  <= "00" & data1(1 downto 0);5�_�  H  J          I   �   *    ����                                                                                                                                                                                                                                                                                                                            �   *       �   -       v   -    ^N   i �   �   �   �      C                        m1_axis_tdata  <= "00" & data1(3 downto 2);�   �   �   �    5�_�  I  K          J   u       ����                                                                                                                                                                                                                                                                                                                            �   *       �   1       v   -    ^�     �   t   v   �    �   u   v   �    5�_�  J  L          K   v       ����                                                                                                                                                                                                                                                                                                                            �   *       �   1       v   -    ^�   j �   u   w   �                  data         := 0;5�_�  K  M          L   }        ����                                                                                                                                                                                                                                                                                                                            }          �          V       ^�     �   |   }          %                     if data2=15 then   #                        data2 := 0;                        else   +                        data2 := data2 + 1;                        end if;5�_�  L  N          M   ~       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   l �   }   �   �    �   ~      �    5�_�  M  O          N   v       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�     �   u   w   �                  data2         := 0;5�_�  N  P          O   v       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   m �   u   w   �                   data2         := 50;5�_�  O  _          P   �   8    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^Y     �   �   �   �      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);5�_�  P  `  Q      _   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^b     �   �   �   �      D                     m1_axis_tdata  <= "000000" & data1(3 downto 0);5�_�  _  a          `   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^c   n �   �   �   �      C                     m1_axis_tdata  <= "00000" & data1(3 downto 0);5�_�  `  b          a   �       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^z     �   �   �   �    �   �   �   �    5�_�  a  c          b   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^|     �   �   �   �      B                     m1_axis_tdata  <= "0000" & data1(3 downto 0);5�_�  b  d          c   �   8    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^     �   �   �   �      D                     m1_axis_tdata  <= "000000" & data1(3 downto 0);5�_�  c  e          d   �       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   p �   �   �   �      B                     m1_axis_tdata  <= "0000" & data1(3 downto 0);5�_�  d  f          e   v       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   q �   u   w   �                  data2         := 5;5�_�  e  g          f   ~       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   r �   }      �      %                     if data2=15 then5�_�  f  h          g   ~       ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^�   s �   }      �      %                     if data2= 4 then5�_�  g  i          h   ~       ����                                                                                                                                                                                                                                                                                                                                                             ^?   t �   }      �      %                     if data2= 3 then5�_�  h  j          i   ~       ����                                                                                                                                                                                                                                                                                                                                                             ^?9   u �   }      �      %                     if data2= 7 then5�_�  i  k          j   ~       ����                                                                                                                                                                                                                                                                                                                                                             ^K�   v �   }      �      %                     if data2= 4 then5�_�  j  l          k   ~       ����                                                                                                                                                                                                                                                                                                                                                             ^L   w �   }      �      %                     if data2= 7 then5�_�  k  m          l   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   �   �   �                   N     => 16,5�_�  l  n          m   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   �   �   �                   N     => 816,5�_�  m  o          n   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   x �   �   �   �                   N     => 86,5�_�  n  p          o   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   �   �   �                   N     => 8,5�_�  o  q          p   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   y �   �   �   �                   N     => 108,5�_�  p  r          q   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   z �   �   �   �                   N     => 10,5�_�  q  s          r   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   { �   �   �   �                   N     => 14,5�_�  r  t          s   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   �   �   �                   N     => 13,5�_�  s  u          t   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   �   �   �                   N     => 1rr5�_�  t  v          u   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   | �   �   �   �                   N     => 12r5�_�  u  w          v   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   } �   �   �   �                   N     => 12,5�_�  v  x          w   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��   ~ �   �   �   �                   N     => 11,5�_�  w  y          x   �       ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   �   �   �                   N     => 12,5�_�  x  z          y   :        ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   9   L   �    �   :   ;   �    5�_�  y  {          z   L        ����                                                                                                                                                                                                                                                                                                                            L           ]          V        ^�     �   \   ^             end component cordic; --}}}�   K   M             component cordic is --{{{5�_�  z  |          {   ^        ����                                                                                                                                                                                                                                                                                                                            L           ]          V        ^�
     �   ]   p   �    �   ^   _   �    5�_�  {  }          |   ^        ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�     �   n   p             end component cordic; --}}}�   ]   _             component cordic is --{{{5�_�  |  ~          }   V   1    ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�      �   U   W   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  }            ~   c   1    ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�(     �   b   d   �      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  ~  �             c   1    ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�T     �   b   d   �      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);5�_�    �          �   h   1    ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�[     �   g   i   �      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            ^           o          V        ^�i     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^�l     �   �   �          cordic_inst:cordic --{{{5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            �           �   4       V        ^�n     �   �        �           5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         4       V        ^�r     �   �            cordic_inst:cordic --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4               ^�     �   �   �            port map(   '           m_axis_tdata  =>axis2_tdata,   (           m_axis_tvalid =>axis2_tvalid,   '           m_axis_tlast  =>axis2_tlast,   (           m_axis_tready =>axis2_tready,   )           s_axis_tdata  =>m1_axis_tdata,   *           s_axis_tvalid =>m1_axis_tvalid,   )           s_axis_tlast  =>m1_axis_tlast,   *           s_axis_tready =>m1_axis_tready,   -           clk           =>clk_tb           ,   4           rst           =>rst_tb           ); --}}}�   �   �        mapper_inst:mapper --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   4               ^��     �   �   �           generic map(                N     => 16,                ITER  => 10)       port map(     '           m_axis_tdata  =>axisO_tdata,   (           m_axis_tvalid =>axisO_tvalid,   '           m_axis_tlast  =>axisO_tlast,   (           m_axis_tready =>axisO_tready,   '           s_axis_tdata  =>axis2_tdata,   (           s_axis_tvalid =>axis2_tvalid,   '           s_axis_tlast  =>axis2_tlast,   (           s_axis_tready =>axis2_tready,   -           clk           =>clk_tb           ,   4           rst           =>rst_tb           ); --}}}�   �   �        cordic_inst:cordic --{{{5�_�  �  �          �   o       ����                                                                                                                                                                                                                                                                                                                            �           �   4               ^��     �   o   q      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^��     �   �   �        (           s_axis_tvalid =>axis2_tvalid,   '           s_axis_tlast  =>axis2_tlast,   (           s_axis_tready =>axis2_tready,�   �   �        '           s_axis_tdata  =>axis2_tdata,5�_�  �  �          �   �   !    ����                                                                                                                                                                                                                                                                                                                            �   !       �   !          !    ^��     �   �   �        )           s_axis_tdata  =>s_axis2_tdata,   *           s_axis_tvalid =>s_axis2_tvalid,   )           s_axis_tlast  =>s_axis2_tlast,   *           s_axis_tready =>s_axis2_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^��     �   �   �        (           s_axis_tdata  =>s_axis_tdata,   )           s_axis_tvalid =>s_axis_tvalid,   (           s_axis_tlast  =>s_axis_tlast,   )           s_axis_tready =>s_axis_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^��     �   �   �        )           s_axis_tvalid =>m_axis_tvalid,   (           s_axis_tlast  =>m_axis_tlast,   )           s_axis_tready =>m_axis_tready,�   �   �        (           s_axis_tdata  =>m_axis_tdata,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^��     �   �   �        '           m_axis_tdata  =>axisO_tdata,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^�   � �   �   �        '           m_axis_tdata  =>axisO_tdata,   (           m_axis_tvalid =>axisO_tvalid,   '           m_axis_tlast  =>axisO_tlast,   (           m_axis_tready =>axisO_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^�X     �   �   �        (           m_axis_tvalid =>axis2_tvalid,   '           m_axis_tlast  =>axis2_tlast,   (           m_axis_tready =>axis2_tready,�   �   �        '           m_axis_tdata  =>axis2_tdata,5�_�  �  �          �   �   !    ����                                                                                                                                                                                                                                                                                                                            �   !       �   !          !    ^�Z     �   �   �        )           m_axis_tdata  =>axis102_tdata,   *           m_axis_tvalid =>axis102_tvalid,   )           m_axis_tlast  =>axis102_tlast,   *           m_axis_tready =>axis102_tready,5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   !       �   !          !    ^�a     �   �   �      �   �   �      5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                                                                                                                            �   !       �   !          !    ^�i     �   �   �        K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  �  �          �   �   ,    ����                                                                                                                                                                                                                                                                                                                            �   !       �   !          !    ^�j     �   �   �        M   signal axis2_tdata:  STD_LOGIC_VECTOR (157 downto 0):=(others=>'0'); --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   -       V       ^�y     �   �   �          -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �          '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �          '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �          L   signal axis2_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   .       V        ^�|     �   �   �      �   �   �      5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �   .       V       ^��     �   �   �          M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{   (   signal axis10_tvalid: STD_LOGIC:='0';   (   signal axis10_tlast:  STD_LOGIC:='0';   .   signal axis10_tready: STD_LOGIC:='0'; --}}}5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     ^��   � �            &           s_axis_tdata  =>axis_tdata,�            '           s_axis_tdata  =>axis2_tdata,   (           s_axis_tvalid =>axis2_tvalid,   '           s_axis_tlast  =>axis2_tlast,   (           s_axis_tready =>axis2_tready,5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                     ^��     �   �   �      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                                                     ^��     �   �   �        --cordic_inst:cordic --{{{5�_�  �  �          �   c   1    ����                                                                                                                                                                                                                                                                                                                                                     ^��   � �   b   d        =           m_axis_tdata  : out STD_LOGIC_VECTOR (8 downto 0);5�_�  �  �  �      �   �        ����                                                                                                                                                                                                                                                                                                                            �                             ^�N   � �   �             generic map(                N     => 16,                ITER  => 10)       port map(     (           m_axis_tdata  =>axis10_tdata,   )           m_axis_tvalid =>axis10_tvalid,   (           m_axis_tlast  =>axis10_tlast,   )           m_axis_tready =>axis10_tready,   )           s_axis_tdata  =>m1_axis_tdata,   *           s_axis_tvalid =>m1_axis_tvalid,   )           s_axis_tlast  =>m1_axis_tlast,   *           s_axis_tready =>m1_axis_tready,   -           clk           =>clk_tb           ,   4           rst           =>rst_tb           ); --}}}�   �   �        $join_16from8_inst:join_16from8 --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �                           ^�[   � �   �          &--join_16from8_inst:join_16from8 --{{{   --   generic map(   --             N     => 16,   --             ITER  => 10)   --    port map(     *--           m_axis_tdata  =>axis10_tdata,   +--           m_axis_tvalid =>axis10_tvalid,   *--           m_axis_tlast  =>axis10_tlast,   +--           m_axis_tready =>axis10_tready,   +--           s_axis_tdata  =>m1_axis_tdata,   ,--           s_axis_tvalid =>m1_axis_tvalid,   +--           s_axis_tlast  =>m1_axis_tlast,   ,--           s_axis_tready =>m1_axis_tready,   /--           clk           =>clk_tb           ,   6--           rst           =>rst_tb           ); --}}}5�_�  �  �          �   V   2    ����                                                                                                                                                                                                                                                                                                                            �                           ^�r   � �   U   W        >           s_axis_tdata  : in  STD_LOGIC_VECTOR (16 downto 0);5�_�  �  �          �   Q   1    ����                                                                                                                                                                                                                                                                                                                            �                           ^��     �   P   R        =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �   V   1    ����                                                                                                                                                                                                                                                                                                                            �                           ^��   � �   U   W        >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^��     �   �   �             generic map(                N     => 16,                ITER  => 10)5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                              V       ^��     �                 generic map(                N     => 16,                ITER  => 10)5�_�  �  �          �   _        ����                                                                                                                                                                                                                                                                                                                            _          a          V       ^��     �   ^   _             generic(   9             N     : natural := 16; --Ancho de la palabra   I             ITER  : natural := 10); -- numero de iteraciones por defecto5�_�  �  �          �   M        ����                                                                                                                                                                                                                                                                                                                            M          O          V       ^��   � �   L   M             generic(   9             N     : natural := 16; --Ancho de la palabra   I             ITER  : natural := 10); -- numero de iteraciones por defecto5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                                                             ^"|     �   Z   \          #   component slice_8from16 is --{{{5�_�  �  �          �   i       ����                                                                                                                                                                                                                                                                                                                                                             ^"|     �   h   j          %   end component slice_8from16; --}}}5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             ^"|     �   �   �          &slice_8from16_inst:slice_8from16 --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             ^"|   � �   �   �          &slice_8from48_inst:slice_8from16 --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                                             ^$.$     �   �   �  
    �   �   �  
    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^$.+     �   �   �        $join_16from8_inst:join_16from8 --{{{5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^$..     �   �   �        $join_16from8_inst:join_48from8 --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^$.J     �   �   �      �   �   �      5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$.M     �   �   �        M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{   (   signal axis10_tvalid: STD_LOGIC:='0';   (   signal axis10_tlast:  STD_LOGIC:='0';   .   signal axis10_tready: STD_LOGIC:='0'; --}}}5�_�  �  �          �   [        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$.l     �   Z   j      �   [   \      5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                            [          [          v       ^$.p     �   Z   \  )      "   component join_16from8 is --{{{5�_�  �  �          �   [       ����                                                                                                                                                                                                                                                                                                                            [          [          v       ^$.t     �   Z   \  )      "   component join_48from8 is --{{{5�_�  �  �          �   ]   1    ����                                                                                                                                                                                                                                                                                                                            ]   1       ]   2       v   2    ^$.~     �   \   ^  )      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);5�_�  �  �          �   ]   2    ����                                                                                                                                                                                                                                                                                                                            ]   1       ]   2       v   2    ^$.�     �   \   ^  )      >           m_axis_tdata  : out STD_LOGIC_VECTOR (48 downto 0);5�_�  �  �          �   b   1    ����                                                                                                                                                                                                                                                                                                                            ]   1       ]   2       v   2    ^$.�     �   a   c  )      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �   q   1    ����                                                                                                                                                                                                                                                                                                                            q   1       q   2       v   2    ^$.�     �   p   r  )      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            q   1       q   2       v   2    ^$.�     �   �   �  )    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            q   1       q   2       v   2    ^$.�     �   �   �  *    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            q   1       q   2       v   2    ^$.�     �   �   �  +    �   �   �  +    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$.�     �   �   �  /      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{   (   signal axis11_tvalid: STD_LOGIC:='0';   (   signal axis11_tlast:  STD_LOGIC:='0';   .   signal axis11_tready: STD_LOGIC:='0'; --}}}5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$.�     �   �   �  /      M   signal axis21_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{   (   signal axis21_tvalid: STD_LOGIC:='0';   (   signal axis21_tlast:  STD_LOGIC:='0';   .   signal axis21_tready: STD_LOGIC:='0'; --}}}5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                                                                                                                            �   +       �   ,       v   ,    ^$.�     �   �   �  /      M   signal axis20_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   +       �   ,       v   ,    ^$.�     �   �   �           5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                                     ^$.�     �      .      (           m_axis_tdata  =>axis10_tdata,   )           m_axis_tvalid =>axis10_tvalid,   (           m_axis_tlast  =>axis10_tlast,   )           m_axis_tready =>axis10_tready,5�_�  �  �  �      �         ����                                                                                                                                                                                                                                                                                                                                       (          (    ^$/     �       .                 s_axis_tdata  =>              s_axis_tvalid =>,              s_axis_tlast  =>              s_axis_tready =>,   -           clk           =>clk_tb           ,�      .    �      .      )           s_axis_tdata  =>m1_axis_tdata,   *           s_axis_tvalid =>m1_axis_tvalid,   )           s_axis_tlast  =>m1_axis_tlast,   *           s_axis_tready =>m1_axis_tready,5�_�  �  �          �  '       ����                                                                                                                                                                                                                                                                                                                           '         *                 ^$/     �  &  +  .      (           s_axis_tdata  =>axis10_tdata,   )           s_axis_tvalid =>axis10_tvalid,   (           s_axis_tlast  =>axis10_tlast,   )           s_axis_tready =>axis10_tready,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &   &          &    ^$/`   � �  "  $  .                 m_axis_tdata  =>�  #  $  .    �  "  '  .      '           m_axis_tdata  =>axisO_tdata,   (           m_axis_tvalid =>axisO_tvalid,   '           m_axis_tlast  =>axisO_tlast,   (           m_axis_tready =>axisO_tready,5�_�  �  �          �   i       ����                                                                                                                                                                                                                                                                                                                            i          i          v       ^$0     �   h   j  .      $   end component join_16from8; --}}}5�_�  �  �          �   i       ����                                                                                                                                                                                                                                                                                                                            i          i          v       ^$0#   � �   h   j  .      $   end component join_48from8; --}}}5�_�  �  �          �  #   (    ����                                                                                                                                                                                                                                                                                                                            i          i          v       ^$06   � �  "  $  .      (           m_axis_tdata  =>s1_axis_tdata5�_�  �  �          �  %   (    ����                                                                                                                                                                                                                                                                                                                            i          i          v       ^$0?   � �  $  &  .      (           m_axis_tlast  =>s1_axis_tdata5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                              v       ^$0g     �      .      %join_16from8_inst:join_48from16 --{{{5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                                              v       ^$0m   � �      .      %join_48from8_inst:join_48from16 --{{{5�_�  �  �          �     (    ����                                                                                                                                                                                                                                                                                                                                              v       ^$0�   � �      .      (           s_axis_tdata  =>axis10_tdata,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$0�   � �  "  '  .      )           m_axis_tdata  =>s1_axis_tdata,   )           m_axis_tvalid =>s1_axis_tdata,   )           m_axis_tlast  =>s1_axis_tdata,   )           m_axis_tready =>s1_axis_tdata,5�_�  �  �  �      �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1;     �  "  '  .      )           m_axis_tdata  =>s0_axis_tdata,   )           m_axis_tvalid =>s0_axis_tdata,   )           m_axis_tlast  =>s0_axis_tdata,   )           m_axis_tready =>s0_axis_tdata,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1>   � �  #  '  .      &           m_axis_tvalid =>axis_tdata,   &           m_axis_tlast  =>axis_tdata,   &           m_axis_tready =>axis_tdata,�  "  $  .      &           m_axis_tdata  =>axis_tdata,5�_�  �  �  �      �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1l     �  "  '  .      '           m_axis_tdata  =>axis0_tdata,   '           m_axis_tvalid =>axis0_tdata,   '           m_axis_tlast  =>axis0_tdata,   '           m_axis_tready =>axis0_tdata,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1n     �  "  $  .      '           m_axis_tdata  =>rxis0_tdata,5�_�  �  �  �      �  '       ����                                                                                                                                                                                                                                                                                                                           '         *   '          '    ^$1y     �  &  +  .      (           s_axis_tdata  =>axis20_tdata,   )           s_axis_tvalid =>axis20_tvalid,   (           s_axis_tlast  =>axis20_tlast,   )           s_axis_tready =>axis20_tready,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &   %          %    ^$1}     �  "  (  .                 m_axis_tdata  =>,              m_axis_tvalid =>,              m_axis_tlast  =>,              m_axis_tready =>,   (           s_axis_tdata  =>axis20_tdata,�  #  $  .    �  "  '  .      '           m_axis_tdata  =>jxis0_tdata,   '           m_axis_tvalid =>rxis0_tdata,   '           m_axis_tlast  =>rxis0_tdata,   '           m_axis_tready =>rxis0_tdata,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &   %          %    ^$1�     �  "  (  .                 m_axis_tdata  =>,              m_axis_tvalid =>,              m_axis_tlast  =>,              m_axis_tready =>,   (           s_axis_tdata  =>axis20_tdata,�  #  $  .    �  "  '  .      '           m_axis_tdata  =>jxis0_tdata,   '           m_axis_tvalid =>rxis0_tdata,   '           m_axis_tlast  =>rxis0_tdata,   '           m_axis_tready =>rxis0_tdata,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�   � �  "  '  .      )           m_axis_tdata  =>axis20_tdata,,   )           m_axis_tvalid =>axis20_tvalid,   )           m_axis_tlast  =>axis20_tlast,,   )           m_axis_tready =>axis20_tready,5�_�  �  �          �  %   &    ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�     �  $  &  .      (           m_axis_tlast  =>axis0_tlast,,5�_�  �  �          �  #   &    ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�   � �  "  $  .      (           m_axis_tdata  =>axis0_tdata,,5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�     �   �    .      )--           m_axis_tlast  =>axisO_tlast,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�     �  "  '  .      '           m_axis_tdata  =>axis0_tdata,   (           m_axis_tvalid =>axis0_tvalid,   '           m_axis_tlast  =>axis0_tlast,   (           m_axis_tready =>axis0_tready,5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$1�   � �  "  '  .      '           m_axis_tdata  =>axisL_tdata,   (           m_axis_tvalid =>axisL_tvalid,   '           m_axis_tlast  =>axisL_tlast,   (           m_axis_tready =>axisL_tready,5�_�  �  �          �   X       ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$21   � �   W   \  .    �   X   Y  .    5�_�  �  �          �  #       ����                                                                                                                                                                                                                                                                                                                            X          Z          V       ^$2I     �  "  &  2    �  #  $  2    5�_�  �  �          �  #        ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2M     �  "  $  5      C           m_axis_config_tdata   out STD_LOGIC_VECTOR (7 downto 0);�  "  &  5      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);   0           m_axis_config_tvalid : out STD_LOGIC;   0           m_axis_config_tready : in  STD_LOGIC;5�_�  �  �          �  #   (    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2b     �  "  $  5      J           m_axis_config_tdata  => '1': out STD_LOGIC_VECTOR (7 downto 0);5�_�  �  �          �  $   '    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2c     �  #  %  5      6           m_axis_config_tvalid => '1': out STD_LOGIC;5�_�  �  �          �  %   &    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2f     �  $  &  5      6           m_axis_config_tready => '1': in  STD_LOGIC;5�_�  �  �  �      �  $   &    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2n     �  #  %  5      '           m_axis_config_tvalid => '1':5�_�  �  �          �  #   &    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2o     �  "  $  5      (           m_axis_config_tdata  => '1': 5�_�  �  �          �  %   &    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2q     �  $  &  5      &           m_axis_config_tready => '1'5�_�  �  �          �  #   #    ����                                                                                                                                                                                                                                                                                                                           #   #      #   %       v   %    ^$2s     �  "  $  5      (           m_axis_config_tdata  => '1', 5�_�  �  �          �  $   $    ����                                                                                                                                                                                                                                                                                                                           #   #      #   %       v   %    ^$2�     �  #  %  5      '           m_axis_config_tvalid => '1',5�_�  �  �          �  $   $    ����                                                                                                                                                                                                                                                                                                                           #   #      #   %       v   %    ^$2�     �  #  %  5      '           m_axis_config_tvalid => '1',5�_�  �  �          �  %   $    ����                                                                                                                                                                                                                                                                                                                           #   #      #   %       v   %    ^$2�   � �  $  &  5      '           m_axis_config_tready => '1',5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                           '   $         $       V   $    ^$2�   � �  2  4  5      4           rst           =>rst_tb           ); --}}}�  1  3  5      -           clk           =>clk_tb           ,�  0  2  5      )           s_axis_tready =>axis20_tready,�  /  1  5      (           s_axis_tlast  =>axis20_tlast,�  .  0  5      )           s_axis_tvalid =>axis20_tvalid,�  -  /  5      (           s_axis_tdata  =>axis20_tdata,�  ,  .  5      (           m_axis_tready =>axisO_tready,�  +  -  5      '           m_axis_tlast  =>axisO_tlast,�  *  ,  5      (           m_axis_tvalid =>axisO_tvalid,�  )  +  5      '           m_axis_tdata  =>axisO_tdata,�  (  *  5          port map(  �  &  (  5      <           rst                  => rst_tb           ); --}}}�  %  '  5      5           clk                  => clk_tb           ,�  $  &  5      '           m_axis_config_tready => '1',�  #  %  5      '           m_axis_config_tvalid => '1',�  "  $  5      .           m_axis_config_tdata  => "00000000",�  !  #  5      1           s_axis_tready        => axis10_tready,�     "  5      0           s_axis_tlast         => axis10_tlast,�    !  5      1           s_axis_tvalid        => axis10_tvalid,�       5      0           s_axis_tdata         => axis10_tdata,�      5      1           m_axis_tready        => axis20_tready,�      5      0           m_axis_tlast         => axis20_tlast,�      5      1           m_axis_tvalid        => axis20_tvalid,�      5      0           m_axis_tdata         => axis20_tdata,�      5          port map(  �      5      4           rst           =>rst_tb           ); --}}}�      5      -           clk           =>clk_tb           ,�      5      *           s_axis_tready =>m1_axis_tready,�      5      )           s_axis_tlast  =>m1_axis_tlast,�      5      *           s_axis_tvalid =>m1_axis_tvalid,�      5      )           s_axis_tdata  =>m1_axis_tdata,�      5      )           m_axis_tready =>axis10_tready,�      5      (           m_axis_tlast  =>axis10_tlast,�      5      )           m_axis_tvalid =>axis10_tvalid,�      5      (           m_axis_tdata  =>axis10_tdata,�      5          port map(  �  
    5      6--           rst           =>rst_tb           ); --}}}�  	    5      /--           clk           =>clk_tb           ,�    
  5      *--           s_axis_tready =>axis2_tready,�    	  5      )--           s_axis_tlast  =>axis2_tlast,�      5      *--           s_axis_tvalid =>axis2_tvalid,�      5      )--           s_axis_tdata  =>axis2_tdata,�      5      *--           m_axis_tready =>axisO_tready,�      5      (--           m_axis_tlast  >axisO_tlast,�      5      *--           m_axis_tvalid =>axisO_tvalid,�      5      )--           m_axis_tdata  =>axisO_tdata,�       5      --    port map(  �   �    5      --             ITER  => 10)�   �     5      --             N     => 16,�   �   �  5      --   generic map(�   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m1_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  5      *--           m_axis_tready =>axis2_tready,�   �   �  5      )--           m_axis_tlast  =>axis2_tlast,�   �   �  5      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  5      )--           m_axis_tdata  =>axis2_tdata,�   �   �  5      --    port map(�   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m3_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  5      ,--           m_axis_tready =>s3_axis_tready,�   �   �  5      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  5      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  5      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  5      --    port map(  �   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m3_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  5      ,--           m_axis_tready =>s3_axis_tready,�   �   �  5      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  5      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  5      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  5      --    port map(  �   �   �  5      %   end process axi_master_proc; --}}}�   �   �  5            end if;�   �   �  5               end if;�   �   �  5                  end case;�   �   �  5                        end if;�   �   �  5                           end if;�   �   �  5      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  5      .                        s1_axis_tready <= '1';�   �   �  5      .                        m1_axis_tvalid <= '0';�   �   �  5                           else�   �   �  5      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  5      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  5      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  5      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  5      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  5      $               when waitingMready =>�   �   �  5                        end if;�   �   �  5      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  5      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  5      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  5      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  5      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  5                           end if;�   �   �  5      +                        data2 := data2 + 1;�   �   �  5                           else�   �   �  5      #                        data2 := 0;�   �   �  5      &                     if data2= 15 then�   �   �  5      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  5      )                     bitCounter     := 0;�   �   �  5      *                     s1_axis_tready <='0';�   �   �  5      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  5      $               when waitingSvalid =>�   �   �  5                  case state is�   �   �  5               else�   �   �  5                  data2         := 0;�   �   �  5                  data         := 0;�   �   �  5      .            m1_axis_tdata  <= (others => '0');�   �   �  5      "            m1_axis_tvalid <= '0';�   �   �  5      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  5      "            s1_axis_tready <= '1';�   �   �  5      ,            state          <= waitingSvalid;�   �   �  5               if rst_tb = '0' then�   �   �  5      !      if rising_edge(clk_tb) then�   �   �  5         begin�   �   �  5      ,      variable data2 :natural range 0 to 15;�   �   �  5      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  5      2      variable data :integer range -128 to 127:=0;�   �   �  5      0      variable bitCounter :integer range 0 to 8;�   �   �  5      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  5          rst_tb   <= '1' after 180 ns;�   �   �  5      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  5      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  5      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  5      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  5      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  5      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  5      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  5      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  5      )   signal m1_axis_tready: STD_LOGIC:='1';�      �  5      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   ~   �  5      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   }     5      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   {   }  5      %   end component slice_8from48; --}}}�   z   |  5      *           rst           : in  STD_LOGIC);�   y   {  5      )           clk           : in  STD_LOGIC;�   w   y  5      )           s_axis_tready : out STD_LOGIC;�   v   x  5      )           s_axis_tlast  : in  STD_LOGIC;�   u   w  5      )           s_axis_tvalid : in  STD_LOGIC;�   t   v  5      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  5      )           m_axis_tready : in  STD_LOGIC;�   q   s  5      )           m_axis_tlast  : out STD_LOGIC;�   p   r  5      )           m_axis_tvalid : out STD_LOGIC;�   o   q  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   n   p  5      	    port(�   m   o  5      #   component slice_8from48 is --{{{�   l   n  5      %   end component join_48from16; --}}}�   k   m  5      *           rst           : in  STD_LOGIC);�   j   l  5      )           clk           : in  STD_LOGIC;�   h   j  5      )           s_axis_tready : out STD_LOGIC;�   g   i  5      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  5      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  5      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (16 downto 0);�   c   e  5      )           m_axis_tready : in  STD_LOGIC;�   b   d  5      )           m_axis_tlast  : out STD_LOGIC;�   a   c  5      )           m_axis_tvalid : out STD_LOGIC;�   `   b  5      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  5      	    port(�   ^   `  5      #   component join_48from16 is --{{{�   ]   _  5      $   end component join_16from8; --}}}�   \   ^  5      *           rst           : in  STD_LOGIC);�   [   ]  5      )           clk           : in  STD_LOGIC;�   Y   [  5      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  5      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  5      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  5      )           s_axis_tready : out STD_LOGIC;�   T   V  5      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  5      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  5      )           m_axis_tready : in  STD_LOGIC;�   O   Q  5      )           m_axis_tlast  : out STD_LOGIC;�   N   P  5      )           m_axis_tvalid : out STD_LOGIC;�   M   O  5      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  5      	    port(�   K   M  5      "   component join_16from8 is --{{{�   J   L  5         end component cordic; --}}}�   I   K  5      *           rst           : in  STD_LOGIC);�   H   J  5      )           clk           : in  STD_LOGIC;�   F   H  5      )           s_axis_tready : out STD_LOGIC;�   E   G  5      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  5      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  5      )           m_axis_tready : in  STD_LOGIC;�   @   B  5      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  5      )           m_axis_tvalid : out STD_LOGIC;�   >   @  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  5      	    port(�   <   >  5      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  5      9             N     : natural := 16; --Ancho de la palabra�   :   <  5         generic(�   9   ;  5         component cordic is --{{{�   8   :  5         end component mapper; --}}}�   7   9  5      *           rst           : in  STD_LOGIC);�   6   8  5      )           clk           : in  STD_LOGIC;�   4   6  5      )           s_axis_tready : out STD_LOGIC;�   3   5  5      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  5      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  5      )           m_axis_tready : in  STD_LOGIC;�   .   0  5      )           m_axis_tlast  : out STD_LOGIC;�   -   /  5      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  5      	    port(�   *   ,  5         component mapper is --{{{�   )   +  5      $   end component slice_2from8; --}}}�   (   *  5      *           rst           : in  STD_LOGIC);�   '   )  5      )           clk           : in  STD_LOGIC;�   %   '  5      )           s_axis_tready : out STD_LOGIC;�   $   &  5      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  5      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  5      )           m_axis_tready : in  STD_LOGIC;�      !  5      )           m_axis_tlast  : out STD_LOGIC;�         5      )           m_axis_tvalid : out STD_LOGIC;�        5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        5      	    port(�        5      "   component slice_2from8 is --{{{�        5      $   end component slice_1from8; --}}}�        5      *           rst           : in  STD_LOGIC);�        5      )           clk           : in  STD_LOGIC;�        5      )           s_axis_tready : out STD_LOGIC;�        5      )           s_axis_tlast  : in  STD_LOGIC;�        5      )           s_axis_tvalid : in  STD_LOGIC;�        5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        5      )           m_axis_tready : in  STD_LOGIC;�        5      )           m_axis_tlast  : out STD_LOGIC;�        5      )           m_axis_tvalid : out STD_LOGIC;�        5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        5      	    port(�        5      "   component slice_1from8 is --{{{�        5      .   signal rst_tb            : STD_LOGIC:= '0';�   
     5      .   signal clk_tb            : STD_LOGIC:= '0';�      
  5      4   signal state   :axiStates := waitingSvalid; --}}}�      	  5      6   type   axiStates is (waitingSvalid, waitingMready);�  !  #          )           s_axis_tready =>axis10_tready,�  "  $          /           m_axis_config_tdata  => "00000000", �  $  &          '           m_axis_config_tready => '1',�              (           m_axis_tlast  =>axis20_tlast,�  %  '          -           clk           =>clk_tb           ,�  #  %          '           m_axis_config_tvalid => '1',�              (           m_axis_tdata  =>axis20_tdata,�              )           m_axis_tvalid =>axis20_tvalid,�  &  (          4           rst           =>rst_tb           ); --}}}�     "          (           s_axis_tlast  =>axis10_tlast,�    !          )           s_axis_tvalid =>axis10_tvalid,�               (           s_axis_tdata  =>axis10_tdata,�              )           m_axis_tready =>axis20_tready,5�_�  �  �          �  #        ����                                                                                                                                                                                                                                                                                                                           #          %           V        ^$2�     �  "  #          .           m_axis_config_tdata  => "00000000",   '           m_axis_config_tvalid => '1',   '           m_axis_config_tready => '1',5�_�  �  �          �         ����                                                                                                                                                                                                                                                                                                                           #          #           V        ^$2�     �      2    �      2    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                              V       ^$2�   � �  2  4  5      4           rst           =>rst_tb           ); --}}}�  1  3  5      -           clk           =>clk_tb           ,�  0  2  5      )           s_axis_tready =>axis20_tready,�  /  1  5      (           s_axis_tlast  =>axis20_tlast,�  .  0  5      )           s_axis_tvalid =>axis20_tvalid,�  -  /  5      (           s_axis_tdata  =>axis20_tdata,�  ,  .  5      (           m_axis_tready =>axisO_tready,�  +  -  5      '           m_axis_tlast  =>axisO_tlast,�  *  ,  5      (           m_axis_tvalid =>axisO_tvalid,�  )  +  5      '           m_axis_tdata  =>axisO_tdata,�  (  *  5          port map(  �  &  (  5      <           rst                  => rst_tb           ); --}}}�  %  '  5      5           clk                  => clk_tb           ,�  $  &  5      1           s_axis_tready        => axis10_tready,�  #  %  5      0           s_axis_tlast         => axis10_tlast,�  "  $  5      1           s_axis_tvalid        => axis10_tvalid,�  !  #  5      0           s_axis_tdata         => axis10_tdata,�     "  5      1           m_axis_tready        => axis20_tready,�    !  5      0           m_axis_tlast         => axis20_tlast,�       5      1           m_axis_tvalid        => axis20_tvalid,�      5      0           m_axis_tdata         => axis20_tdata,�      5          port map(  �      5      <           rst                  => rst_tb           ); --}}}�      5      5           clk                  => clk_tb           ,�      5      '           m_axis_config_tready => '1',�      5      '           m_axis_config_tvalid => '1',�      5      .           m_axis_config_tdata  => "00000000",�      5      2           s_axis_tready        => m1_axis_tready,�      5      1           s_axis_tlast         => m1_axis_tlast,�      5      2           s_axis_tvalid        => m1_axis_tvalid,�      5      1           s_axis_tdata         => m1_axis_tdata,�      5      1           m_axis_tready        => axis10_tready,�      5      0           m_axis_tlast         => axis10_tlast,�      5      1           m_axis_tvalid        => axis10_tvalid,�      5      0           m_axis_tdata         => axis10_tdata,�      5          port map(  �  
    5      6--           rst           =>rst_tb           ); --}}}�  	    5      /--           clk           =>clk_tb           ,�    
  5      *--           s_axis_tready =>axis2_tready,�    	  5      )--           s_axis_tlast  =>axis2_tlast,�      5      *--           s_axis_tvalid =>axis2_tvalid,�      5      )--           s_axis_tdata  =>axis2_tdata,�      5      *--           m_axis_tready =>axisO_tready,�      5      (--           m_axis_tlast  >axisO_tlast,�      5      *--           m_axis_tvalid =>axisO_tvalid,�      5      )--           m_axis_tdata  =>axisO_tdata,�       5      --    port map(  �   �    5      --             ITER  => 10)�   �     5      --             N     => 16,�   �   �  5      --   generic map(�   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m1_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  5      *--           m_axis_tready =>axis2_tready,�   �   �  5      )--           m_axis_tlast  =>axis2_tlast,�   �   �  5      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  5      )--           m_axis_tdata  =>axis2_tdata,�   �   �  5      --    port map(�   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m3_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  5      ,--           m_axis_tready =>s3_axis_tready,�   �   �  5      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  5      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  5      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  5      --    port map(  �   �   �  5      6--           rst           =>rst_tb           ); --}}}�   �   �  5      /--           clk           =>clk_tb           ,�   �   �  5      ,--           s_axis_tready =>m3_axis_tready,�   �   �  5      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  5      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  5      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  5      ,--           m_axis_tready =>s3_axis_tready,�   �   �  5      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  5      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  5      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  5      --    port map(  �   �   �  5      %   end process axi_master_proc; --}}}�   �   �  5            end if;�   �   �  5               end if;�   �   �  5                  end case;�   �   �  5                        end if;�   �   �  5                           end if;�   �   �  5      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  5      .                        s1_axis_tready <= '1';�   �   �  5      .                        m1_axis_tvalid <= '0';�   �   �  5                           else�   �   �  5      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  5      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  5      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  5      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  5      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  5      $               when waitingMready =>�   �   �  5                        end if;�   �   �  5      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  5      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  5      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  5      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  5      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  5                           end if;�   �   �  5      +                        data2 := data2 + 1;�   �   �  5                           else�   �   �  5      #                        data2 := 0;�   �   �  5      &                     if data2= 15 then�   �   �  5      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  5      )                     bitCounter     := 0;�   �   �  5      *                     s1_axis_tready <='0';�   �   �  5      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  5      $               when waitingSvalid =>�   �   �  5                  case state is�   �   �  5               else�   �   �  5                  data2         := 0;�   �   �  5                  data         := 0;�   �   �  5      .            m1_axis_tdata  <= (others => '0');�   �   �  5      "            m1_axis_tvalid <= '0';�   �   �  5      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  5      "            s1_axis_tready <= '1';�   �   �  5      ,            state          <= waitingSvalid;�   �   �  5               if rst_tb = '0' then�   �   �  5      !      if rising_edge(clk_tb) then�   �   �  5         begin�   �   �  5      ,      variable data2 :natural range 0 to 15;�   �   �  5      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  5      2      variable data :integer range -128 to 127:=0;�   �   �  5      0      variable bitCounter :integer range 0 to 8;�   �   �  5      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  5          rst_tb   <= '1' after 180 ns;�   �   �  5      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  5      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  5      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  5      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  5      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  5      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  5      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  5      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  5      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  5      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  5      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  5      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  5      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  5      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  5      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  5      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  5      )   signal m1_axis_tready: STD_LOGIC:='1';�      �  5      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   ~   �  5      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   }     5      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   {   }  5      %   end component slice_8from48; --}}}�   z   |  5      *           rst           : in  STD_LOGIC);�   y   {  5      )           clk           : in  STD_LOGIC;�   w   y  5      )           s_axis_tready : out STD_LOGIC;�   v   x  5      )           s_axis_tlast  : in  STD_LOGIC;�   u   w  5      )           s_axis_tvalid : in  STD_LOGIC;�   t   v  5      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  5      )           m_axis_tready : in  STD_LOGIC;�   q   s  5      )           m_axis_tlast  : out STD_LOGIC;�   p   r  5      )           m_axis_tvalid : out STD_LOGIC;�   o   q  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   n   p  5      	    port(�   m   o  5      #   component slice_8from48 is --{{{�   l   n  5      %   end component join_48from16; --}}}�   k   m  5      *           rst           : in  STD_LOGIC);�   j   l  5      )           clk           : in  STD_LOGIC;�   h   j  5      )           s_axis_tready : out STD_LOGIC;�   g   i  5      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  5      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  5      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (16 downto 0);�   c   e  5      )           m_axis_tready : in  STD_LOGIC;�   b   d  5      )           m_axis_tlast  : out STD_LOGIC;�   a   c  5      )           m_axis_tvalid : out STD_LOGIC;�   `   b  5      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  5      	    port(�   ^   `  5      #   component join_48from16 is --{{{�   ]   _  5      $   end component join_16from8; --}}}�   \   ^  5      *           rst           : in  STD_LOGIC);�   [   ]  5      )           clk           : in  STD_LOGIC;�   Y   [  5      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  5      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  5      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  5      )           s_axis_tready : out STD_LOGIC;�   T   V  5      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  5      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  5      )           m_axis_tready : in  STD_LOGIC;�   O   Q  5      )           m_axis_tlast  : out STD_LOGIC;�   N   P  5      )           m_axis_tvalid : out STD_LOGIC;�   M   O  5      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  5      	    port(�   K   M  5      "   component join_16from8 is --{{{�   J   L  5         end component cordic; --}}}�   I   K  5      *           rst           : in  STD_LOGIC);�   H   J  5      )           clk           : in  STD_LOGIC;�   F   H  5      )           s_axis_tready : out STD_LOGIC;�   E   G  5      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  5      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  5      )           m_axis_tready : in  STD_LOGIC;�   @   B  5      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  5      )           m_axis_tvalid : out STD_LOGIC;�   >   @  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  5      	    port(�   <   >  5      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  5      9             N     : natural := 16; --Ancho de la palabra�   :   <  5         generic(�   9   ;  5         component cordic is --{{{�   8   :  5         end component mapper; --}}}�   7   9  5      *           rst           : in  STD_LOGIC);�   6   8  5      )           clk           : in  STD_LOGIC;�   4   6  5      )           s_axis_tready : out STD_LOGIC;�   3   5  5      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  5      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  5      )           m_axis_tready : in  STD_LOGIC;�   .   0  5      )           m_axis_tlast  : out STD_LOGIC;�   -   /  5      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  5      	    port(�   *   ,  5         component mapper is --{{{�   )   +  5      $   end component slice_2from8; --}}}�   (   *  5      *           rst           : in  STD_LOGIC);�   '   )  5      )           clk           : in  STD_LOGIC;�   %   '  5      )           s_axis_tready : out STD_LOGIC;�   $   &  5      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  5      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  5      )           m_axis_tready : in  STD_LOGIC;�      !  5      )           m_axis_tlast  : out STD_LOGIC;�         5      )           m_axis_tvalid : out STD_LOGIC;�        5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        5      	    port(�        5      "   component slice_2from8 is --{{{�        5      $   end component slice_1from8; --}}}�        5      *           rst           : in  STD_LOGIC);�        5      )           clk           : in  STD_LOGIC;�        5      )           s_axis_tready : out STD_LOGIC;�        5      )           s_axis_tlast  : in  STD_LOGIC;�        5      )           s_axis_tvalid : in  STD_LOGIC;�        5      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        5      )           m_axis_tready : in  STD_LOGIC;�        5      )           m_axis_tlast  : out STD_LOGIC;�        5      )           m_axis_tvalid : out STD_LOGIC;�        5      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        5      	    port(�        5      "   component slice_1from8 is --{{{�        5      .   signal rst_tb            : STD_LOGIC:= '0';�   
     5      .   signal clk_tb            : STD_LOGIC:= '0';�      
  5      4   signal state   :axiStates := waitingSvalid; --}}}�      	  5      6   type   axiStates is (waitingSvalid, waitingMready);�              *           s_axis_tready =>m1_axis_tready,�              .           m_axis_config_tdata  => "00000000",�              )           s_axis_tdata  =>m1_axis_tdata,�              -           clk           =>clk_tb           ,�              '           m_axis_config_tready => '1',�              '           m_axis_config_tvalid => '1',�              )           m_axis_tready =>axis10_tready,�              (           m_axis_tlast  =>axis10_tlast,�              )           m_axis_tvalid =>axis10_tvalid,�              (           m_axis_tdata  =>axis10_tdata,�              *           s_axis_tvalid =>m1_axis_tvalid,�              4           rst           =>rst_tb           ); --}}}�              )           s_axis_tlast  =>m1_axis_tlast,5�_�  �  �  �      �     #    ����                                                                                                                                                                                                                                                                                                                              #         -       v   -    ^$B�     �      5      .           m_axis_config_tdata  => "00000000",�      5    5�_�  �  �          �     /    ����                                                                                                                                                                                                                                                                                                                              #         .       v   -    ^$B�     �      5      /           m_axis_config_tdata  => axis10_tdata5�_�  �  �          �     (    ����                                                                                                                                                                                                                                                                                                                              #         .       v   -    ^$B�     �      5      0           m_axis_config_tdata  => axis10_tdata,5�_�  �  �          �     #    ����                                                                                                                                                                                                                                                                                                                              #         %       v   %    ^$B�     �      5      '           m_axis_config_tvalid => '1',�      5    5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                              +         .       v   .    ^$B�     �      5      0           m_axis_config_tvalid => axis11_tdata,5�_�  �  �          �     #    ����                                                                                                                                                                                                                                                                                                                              #         %       v   %    ^$B�     �      5      '           m_axis_config_tready => '1',�      5    5�_�  �  �          �     +    ����                                                                                                                                                                                                                                                                                                                              #         /       v   %    ^$B�   � �      5      1           m_axis_config_tready => axis11_tvalid,5�_�  �  �          �     '    ����                                                                                                                                                                                                                                                                                                                              '         '          '    ^$B�     �      5      /           m_axis_config_tdata  => axis1_tdata,�      5      0           m_axis_config_tdata  => axis11_tdata,   1           m_axis_config_tvalid => axis11_tvalid,   1           m_axis_config_tready => axis11_tready,5�_�  �  �          �     (    ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$B�   � �      5      0           m_axis_config_tdata  => axis41_tdata,   1           m_axis_config_tvalid => axis41_tvalid,   1           m_axis_config_tready => axis41_tready,5�_�  �  �          �   f   2    ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$B�   � �   e   g  5      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (16 downto 0);5�_�  �  �  �      �  2        ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$Cy     �  1  5  5    �  2  3  5    5�_�  �  �          �  2        ����                                                                                                                                                                                                                                                                                                                           2          4   $          $    ^$C|     �  1  3  8      ?           m_axis_config_tdata   STD_LOGIC_VECTOR (7 downto 0);�  1  5  8      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);   0           m_axis_config_tvalid : out STD_LOGIC;   0           m_axis_config_tready : in  STD_LOGIC;5�_�  �  �          �  2   #    ����                                                                                                                                                                                                                                                                                                                           2   #      4   #          #    ^$C�     �  2  5  8      -           m_axis_config_tvalid => STD_LOGIC;   -           m_axis_config_tready => STD_LOGIC;�  1  3  8      A           m_axis_config_tdata  => STD_LOGIC_VECTOR (7 downto 0);5�_�  �             �  2   .    ����                                                                                                                                                                                                                                                                                                                           2   #      4   #          #    ^$C�     �  1  3  8      L           m_axis_config_tdata  => axis3_tdataSTD_LOGIC_VECTOR (7 downto 0);5�_�  �               3   .    ����                                                                                                                                                                                                                                                                                                                           2   #      4   #          #    ^$C�     �  2  4  8      8           m_axis_config_tvalid => axis3_tdataSTD_LOGIC;5�_�                 4   .    ����                                                                                                                                                                                                                                                                                                                           2   #      4   #          #    ^$C�     �  3  5  8      8           m_axis_config_tready => axis3_tdataSTD_LOGIC;5�_�                2   .    ����                                                                                                                                                                                                                                                                                                                           2   .      4   .          .    ^$C�     �  1  5  8      /           m_axis_config_tdata  => axis3_tdata;   /           m_axis_config_tvalid => axis3_tdata;   /           m_axis_config_tready => axis3_tdata;5�_�                3   *    ����                                                                                                                                                                                                                                                                                                                           2   .      4   .          .    ^$C�     �  2  4  8      /           m_axis_config_tvalid => axis3_tdata,5�_�                4   *    ����                                                                                                                                                                                                                                                                                                                           2   .      4   .          .    ^$C�   � �  3  5  8      /           m_axis_config_tready => axis3_tdata,5�_�                *        ����                                                                                                                                                                                                                                                                                                                           6   .      *          V       ^$C�   � �  5  7  8      <           rst                  => rst_tb           ); --}}}�  4  6  8      5           clk                  => clk_tb           ,�  3  5  8      0           m_axis_config_tready => axis3_tready,�  2  4  8      0           m_axis_config_tvalid => axis3_tvalid,�  1  3  8      /           m_axis_config_tdata  => axis3_tdata,�  0  2  8      1           s_axis_tready        => axis20_tready,�  /  1  8      0           s_axis_tlast         => axis20_tlast,�  .  0  8      1           s_axis_tvalid        => axis20_tvalid,�  -  /  8      0           s_axis_tdata         => axis20_tdata,�  ,  .  8      0           m_axis_tready        => axisO_tready,�  +  -  8      /           m_axis_tlast         => axisO_tlast,�  *  ,  8      0           m_axis_tvalid        => axisO_tvalid,�  )  +  8      /           m_axis_tdata         => axisO_tdata,�  (  *  8          port map(  �  &  (  8      <           rst                  => rst_tb           ); --}}}�  %  '  8      5           clk                  => clk_tb           ,�  $  &  8      1           s_axis_tready        => axis10_tready,�  #  %  8      0           s_axis_tlast         => axis10_tlast,�  "  $  8      1           s_axis_tvalid        => axis10_tvalid,�  !  #  8      0           s_axis_tdata         => axis10_tdata,�     "  8      1           m_axis_tready        => axis20_tready,�    !  8      0           m_axis_tlast         => axis20_tlast,�       8      1           m_axis_tvalid        => axis20_tvalid,�      8      0           m_axis_tdata         => axis20_tdata,�      8          port map(  �      8      <           rst                  => rst_tb           ); --}}}�      8      5           clk                  => clk_tb           ,�      8      0           m_axis_config_tready => axis4_tready,�      8      0           m_axis_config_tvalid => axis4_tvalid,�      8      /           m_axis_config_tdata  => axis4_tdata,�      8      2           s_axis_tready        => m1_axis_tready,�      8      1           s_axis_tlast         => m1_axis_tlast,�      8      2           s_axis_tvalid        => m1_axis_tvalid,�      8      1           s_axis_tdata         => m1_axis_tdata,�      8      1           m_axis_tready        => axis10_tready,�      8      0           m_axis_tlast         => axis10_tlast,�      8      1           m_axis_tvalid        => axis10_tvalid,�      8      0           m_axis_tdata         => axis10_tdata,�      8          port map(  �  
    8      6--           rst           =>rst_tb           ); --}}}�  	    8      /--           clk           =>clk_tb           ,�    
  8      *--           s_axis_tready =>axis2_tready,�    	  8      )--           s_axis_tlast  =>axis2_tlast,�      8      *--           s_axis_tvalid =>axis2_tvalid,�      8      )--           s_axis_tdata  =>axis2_tdata,�      8      *--           m_axis_tready =>axisO_tready,�      8      (--           m_axis_tlast  >axisO_tlast,�      8      *--           m_axis_tvalid =>axisO_tvalid,�      8      )--           m_axis_tdata  =>axisO_tdata,�       8      --    port map(  �   �    8      --             ITER  => 10)�   �     8      --             N     => 16,�   �   �  8      --   generic map(�   �   �  8      6--           rst           =>rst_tb           ); --}}}�   �   �  8      /--           clk           =>clk_tb           ,�   �   �  8      ,--           s_axis_tready =>m1_axis_tready,�   �   �  8      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  8      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  8      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  8      *--           m_axis_tready =>axis2_tready,�   �   �  8      )--           m_axis_tlast  =>axis2_tlast,�   �   �  8      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  8      )--           m_axis_tdata  =>axis2_tdata,�   �   �  8      --    port map(�   �   �  8      6--           rst           =>rst_tb           ); --}}}�   �   �  8      /--           clk           =>clk_tb           ,�   �   �  8      ,--           s_axis_tready =>m3_axis_tready,�   �   �  8      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  8      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  8      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  8      ,--           m_axis_tready =>s3_axis_tready,�   �   �  8      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  8      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  8      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  8      --    port map(  �   �   �  8      6--           rst           =>rst_tb           ); --}}}�   �   �  8      /--           clk           =>clk_tb           ,�   �   �  8      ,--           s_axis_tready =>m3_axis_tready,�   �   �  8      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  8      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  8      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  8      ,--           m_axis_tready =>s3_axis_tready,�   �   �  8      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  8      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  8      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  8      --    port map(  �   �   �  8      %   end process axi_master_proc; --}}}�   �   �  8            end if;�   �   �  8               end if;�   �   �  8                  end case;�   �   �  8                        end if;�   �   �  8                           end if;�   �   �  8      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  8      .                        s1_axis_tready <= '1';�   �   �  8      .                        m1_axis_tvalid <= '0';�   �   �  8                           else�   �   �  8      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  8      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  8      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  8      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  8      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  8      $               when waitingMready =>�   �   �  8                        end if;�   �   �  8      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  8      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  8      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  8      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  8      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  8                           end if;�   �   �  8      +                        data2 := data2 + 1;�   �   �  8                           else�   �   �  8      #                        data2 := 0;�   �   �  8      &                     if data2= 15 then�   �   �  8      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  8      )                     bitCounter     := 0;�   �   �  8      *                     s1_axis_tready <='0';�   �   �  8      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  8      $               when waitingSvalid =>�   �   �  8                  case state is�   �   �  8               else�   �   �  8                  data2         := 0;�   �   �  8                  data         := 0;�   �   �  8      .            m1_axis_tdata  <= (others => '0');�   �   �  8      "            m1_axis_tvalid <= '0';�   �   �  8      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  8      "            s1_axis_tready <= '1';�   �   �  8      ,            state          <= waitingSvalid;�   �   �  8               if rst_tb = '0' then�   �   �  8      !      if rising_edge(clk_tb) then�   �   �  8         begin�   �   �  8      ,      variable data2 :natural range 0 to 15;�   �   �  8      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  8      2      variable data :integer range -128 to 127:=0;�   �   �  8      0      variable bitCounter :integer range 0 to 8;�   �   �  8      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  8          rst_tb   <= '1' after 180 ns;�   �   �  8      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  8      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  8      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  8      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  8      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  8      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  8      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  8      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  8      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  8      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  8      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  8      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  8      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  8      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  8      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  8      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  8      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  8      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  8      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  8      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  8      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  8      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  8      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  8      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  8      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  8      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  8      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  8      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  8      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  8      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  8      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  8      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  8      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  8      )   signal m1_axis_tready: STD_LOGIC:='1';�      �  8      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   ~   �  8      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   }     8      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   {   }  8      %   end component slice_8from48; --}}}�   z   |  8      *           rst           : in  STD_LOGIC);�   y   {  8      )           clk           : in  STD_LOGIC;�   w   y  8      )           s_axis_tready : out STD_LOGIC;�   v   x  8      )           s_axis_tlast  : in  STD_LOGIC;�   u   w  8      )           s_axis_tvalid : in  STD_LOGIC;�   t   v  8      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  8      )           m_axis_tready : in  STD_LOGIC;�   q   s  8      )           m_axis_tlast  : out STD_LOGIC;�   p   r  8      )           m_axis_tvalid : out STD_LOGIC;�   o   q  8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   n   p  8      	    port(�   m   o  8      #   component slice_8from48 is --{{{�   l   n  8      %   end component join_48from16; --}}}�   k   m  8      *           rst           : in  STD_LOGIC);�   j   l  8      )           clk           : in  STD_LOGIC;�   h   j  8      )           s_axis_tready : out STD_LOGIC;�   g   i  8      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  8      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  8      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  8      )           m_axis_tready : in  STD_LOGIC;�   b   d  8      )           m_axis_tlast  : out STD_LOGIC;�   a   c  8      )           m_axis_tvalid : out STD_LOGIC;�   `   b  8      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  8      	    port(�   ^   `  8      #   component join_48from16 is --{{{�   ]   _  8      $   end component join_16from8; --}}}�   \   ^  8      *           rst           : in  STD_LOGIC);�   [   ]  8      )           clk           : in  STD_LOGIC;�   Y   [  8      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  8      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  8      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  8      )           s_axis_tready : out STD_LOGIC;�   T   V  8      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  8      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  8      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  8      )           m_axis_tready : in  STD_LOGIC;�   O   Q  8      )           m_axis_tlast  : out STD_LOGIC;�   N   P  8      )           m_axis_tvalid : out STD_LOGIC;�   M   O  8      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  8      	    port(�   K   M  8      "   component join_16from8 is --{{{�   J   L  8         end component cordic; --}}}�   I   K  8      *           rst           : in  STD_LOGIC);�   H   J  8      )           clk           : in  STD_LOGIC;�   F   H  8      )           s_axis_tready : out STD_LOGIC;�   E   G  8      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  8      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  8      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  8      )           m_axis_tready : in  STD_LOGIC;�   @   B  8      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  8      )           m_axis_tvalid : out STD_LOGIC;�   >   @  8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  8      	    port(�   <   >  8      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  8      9             N     : natural := 16; --Ancho de la palabra�   :   <  8         generic(�   9   ;  8         component cordic is --{{{�   8   :  8         end component mapper; --}}}�   7   9  8      *           rst           : in  STD_LOGIC);�   6   8  8      )           clk           : in  STD_LOGIC;�   4   6  8      )           s_axis_tready : out STD_LOGIC;�   3   5  8      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  8      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  8      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  8      )           m_axis_tready : in  STD_LOGIC;�   .   0  8      )           m_axis_tlast  : out STD_LOGIC;�   -   /  8      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  8      	    port(�   *   ,  8         component mapper is --{{{�   )   +  8      $   end component slice_2from8; --}}}�   (   *  8      *           rst           : in  STD_LOGIC);�   '   )  8      )           clk           : in  STD_LOGIC;�   %   '  8      )           s_axis_tready : out STD_LOGIC;�   $   &  8      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  8      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  8      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  8      )           m_axis_tready : in  STD_LOGIC;�      !  8      )           m_axis_tlast  : out STD_LOGIC;�         8      )           m_axis_tvalid : out STD_LOGIC;�        8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        8      	    port(�        8      "   component slice_2from8 is --{{{�        8      $   end component slice_1from8; --}}}�        8      *           rst           : in  STD_LOGIC);�        8      )           clk           : in  STD_LOGIC;�        8      )           s_axis_tready : out STD_LOGIC;�        8      )           s_axis_tlast  : in  STD_LOGIC;�        8      )           s_axis_tvalid : in  STD_LOGIC;�        8      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        8      )           m_axis_tready : in  STD_LOGIC;�        8      )           m_axis_tlast  : out STD_LOGIC;�        8      )           m_axis_tvalid : out STD_LOGIC;�        8      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        8      	    port(�        8      "   component slice_1from8 is --{{{�        8      .   signal rst_tb            : STD_LOGIC:= '0';�   
     8      .   signal clk_tb            : STD_LOGIC:= '0';�      
  8      4   signal state   :axiStates := waitingSvalid; --}}}�      	  8      6   type   axiStates is (waitingSvalid, waitingMready);�  /  1          (           s_axis_tlast  =>axis20_tlast,�  .  0          )           s_axis_tvalid =>axis20_tvalid,�  -  /          (           s_axis_tdata  =>axis20_tdata,�  ,  .          (           m_axis_tready =>axisO_tready,�  +  -          '           m_axis_tlast  =>axisO_tlast,�  *  ,          (           m_axis_tvalid =>axisO_tvalid,�  )  +          '           m_axis_tdata  =>axisO_tdata,�  5  7          4           rst           =>rst_tb           ); --}}}�  4  6          -           clk           =>clk_tb           ,�  3  5          0           m_axis_config_tready => axis3_tready,�  2  4          0           m_axis_config_tvalid => axis3_tvalid,�  1  3          /           m_axis_config_tdata  => axis3_tdata,�  0  2          )           s_axis_tready =>axis20_tready,5�_�                 z       ����                                                                                                                                                                                                                                                                                                                           6   .      *          V       ^$C�     �   y   }  8    �   z   {  8    5�_�                 |       ����                                                                                                                                                                                                                                                                                                                           9   .      -          V       ^$C�     �   |   ~  ;    5�_�    	             p       ����                                                                                                                                                                                                                                                                                                                            p          p          v       ^$C�     �   o   q  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�              	   p        ����                                                                                                                                                                                                                                                                                                                            p                    V       ^$C�   � �  9  ;  <      <           rst                  => rst_tb           ); --}}}�  8  :  <      5           clk                  => clk_tb           ,�  7  9  <      0           m_axis_config_tready => axis3_tready,�  6  8  <      0           m_axis_config_tvalid => axis3_tvalid,�  5  7  <      /           m_axis_config_tdata  => axis3_tdata,�  4  6  <      1           s_axis_tready        => axis20_tready,�  3  5  <      0           s_axis_tlast         => axis20_tlast,�  2  4  <      1           s_axis_tvalid        => axis20_tvalid,�  1  3  <      0           s_axis_tdata         => axis20_tdata,�  0  2  <      0           m_axis_tready        => axisO_tready,�  /  1  <      /           m_axis_tlast         => axisO_tlast,�  .  0  <      0           m_axis_tvalid        => axisO_tvalid,�  -  /  <      /           m_axis_tdata         => axisO_tdata,�  ,  .  <          port map(  �  *  ,  <      <           rst                  => rst_tb           ); --}}}�  )  +  <      5           clk                  => clk_tb           ,�  (  *  <      1           s_axis_tready        => axis10_tready,�  '  )  <      0           s_axis_tlast         => axis10_tlast,�  &  (  <      1           s_axis_tvalid        => axis10_tvalid,�  %  '  <      0           s_axis_tdata         => axis10_tdata,�  $  &  <      1           m_axis_tready        => axis20_tready,�  #  %  <      0           m_axis_tlast         => axis20_tlast,�  "  $  <      1           m_axis_tvalid        => axis20_tvalid,�  !  #  <      0           m_axis_tdata         => axis20_tdata,�     "  <          port map(  �       <      <           rst                  => rst_tb           ); --}}}�      <      5           clk                  => clk_tb           ,�      <      0           m_axis_config_tready => axis4_tready,�      <      0           m_axis_config_tvalid => axis4_tvalid,�      <      /           m_axis_config_tdata  => axis4_tdata,�      <      2           s_axis_tready        => m1_axis_tready,�      <      1           s_axis_tlast         => m1_axis_tlast,�      <      2           s_axis_tvalid        => m1_axis_tvalid,�      <      1           s_axis_tdata         => m1_axis_tdata,�      <      1           m_axis_tready        => axis10_tready,�      <      0           m_axis_tlast         => axis10_tlast,�      <      1           m_axis_tvalid        => axis10_tvalid,�      <      0           m_axis_tdata         => axis10_tdata,�      <          port map(  �      <      6--           rst           =>rst_tb           ); --}}}�      <      /--           clk           =>clk_tb           ,�      <      *--           s_axis_tready =>axis2_tready,�      <      )--           s_axis_tlast  =>axis2_tlast,�  
    <      *--           s_axis_tvalid =>axis2_tvalid,�  	    <      )--           s_axis_tdata  =>axis2_tdata,�    
  <      *--           m_axis_tready =>axisO_tready,�    	  <      (--           m_axis_tlast  >axisO_tlast,�      <      *--           m_axis_tvalid =>axisO_tvalid,�      <      )--           m_axis_tdata  =>axisO_tdata,�      <      --    port map(  �      <      --             ITER  => 10)�      <      --             N     => 16,�      <      --   generic map(�   �    <      6--           rst           =>rst_tb           ); --}}}�   �     <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m1_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  <      *--           m_axis_tready =>axis2_tready,�   �   �  <      )--           m_axis_tlast  =>axis2_tlast,�   �   �  <      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  <      )--           m_axis_tdata  =>axis2_tdata,�   �   �  <      --    port map(�   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      %   end process axi_master_proc; --}}}�   �   �  <            end if;�   �   �  <               end if;�   �   �  <                  end case;�   �   �  <                        end if;�   �   �  <                           end if;�   �   �  <      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      .                        s1_axis_tready <= '1';�   �   �  <      .                        m1_axis_tvalid <= '0';�   �   �  <                           else�   �   �  <      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  <      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  <      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  <      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  <      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  <      $               when waitingMready =>�   �   �  <                        end if;�   �   �  <      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  <      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  <      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  <      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  <                           end if;�   �   �  <      +                        data2 := data2 + 1;�   �   �  <                           else�   �   �  <      #                        data2 := 0;�   �   �  <      &                     if data2= 15 then�   �   �  <      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  <      )                     bitCounter     := 0;�   �   �  <      *                     s1_axis_tready <='0';�   �   �  <      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  <      $               when waitingSvalid =>�   �   �  <                  case state is�   �   �  <               else�   �   �  <                  data2         := 0;�   �   �  <                  data         := 0;�   �   �  <      .            m1_axis_tdata  <= (others => '0');�   �   �  <      "            m1_axis_tvalid <= '0';�   �   �  <      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  <      "            s1_axis_tready <= '1';�   �   �  <      ,            state          <= waitingSvalid;�   �   �  <               if rst_tb = '0' then�   �   �  <      !      if rising_edge(clk_tb) then�   �   �  <         begin�   �   �  <      ,      variable data2 :natural range 0 to 15;�   �   �  <      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  <      2      variable data :integer range -128 to 127:=0;�   �   �  <      0      variable bitCounter :integer range 0 to 8;�   �   �  <      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  <          rst_tb   <= '1' after 180 ns;�   �   �  <      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  <      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  <      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  <      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  <      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  <      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  <      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  <      )   signal m1_axis_tready: STD_LOGIC:='1';�   �   �  <      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�      �  <      %   end component slice_8from48; --}}}�   ~   �  <      1           rst                  : in  STD_LOGIC);�   }     <      0           clk                  : in  STD_LOGIC;�   {   }  <      0           m_axis_config_tready : in  STD_LOGIC;�   z   |  <      0           m_axis_config_tvalid : out STD_LOGIC;�   y   {  <      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�   w   y  <      0           s_axis_tready        : out STD_LOGIC;�   v   x  <      0           s_axis_tlast         : in  STD_LOGIC;�   u   w  <      0           s_axis_tvalid        : in  STD_LOGIC;�   t   v  <      E           s_axis_tdata         : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  <      0           m_axis_tready        : in  STD_LOGIC;�   q   s  <      0           m_axis_tlast         : out STD_LOGIC;�   p   r  <      0           m_axis_tvalid        : out STD_LOGIC;�   o   q  <      E           e_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);�   n   p  <      	    port(�   m   o  <      #   component slice_8from48 is --{{{�   l   n  <      %   end component join_48from16; --}}}�   k   m  <      *           rst           : in  STD_LOGIC);�   j   l  <      )           clk           : in  STD_LOGIC;�   h   j  <      )           s_axis_tready : out STD_LOGIC;�   g   i  <      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  <      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  <      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  <      )           m_axis_tready : in  STD_LOGIC;�   b   d  <      )           m_axis_tlast  : out STD_LOGIC;�   a   c  <      )           m_axis_tvalid : out STD_LOGIC;�   `   b  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  <      	    port(�   ^   `  <      #   component join_48from16 is --{{{�   ]   _  <      $   end component join_16from8; --}}}�   \   ^  <      *           rst           : in  STD_LOGIC);�   [   ]  <      )           clk           : in  STD_LOGIC;�   Y   [  <      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  <      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  <      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  <      )           s_axis_tready : out STD_LOGIC;�   T   V  <      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  <      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  <      )           m_axis_tready : in  STD_LOGIC;�   O   Q  <      )           m_axis_tlast  : out STD_LOGIC;�   N   P  <      )           m_axis_tvalid : out STD_LOGIC;�   M   O  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  <      	    port(�   K   M  <      "   component join_16from8 is --{{{�   J   L  <         end component cordic; --}}}�   I   K  <      *           rst           : in  STD_LOGIC);�   H   J  <      )           clk           : in  STD_LOGIC;�   F   H  <      )           s_axis_tready : out STD_LOGIC;�   E   G  <      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  <      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  <      )           m_axis_tready : in  STD_LOGIC;�   @   B  <      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  <      )           m_axis_tvalid : out STD_LOGIC;�   >   @  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  <      	    port(�   <   >  <      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  <      9             N     : natural := 16; --Ancho de la palabra�   :   <  <         generic(�   9   ;  <         component cordic is --{{{�   8   :  <         end component mapper; --}}}�   7   9  <      *           rst           : in  STD_LOGIC);�   6   8  <      )           clk           : in  STD_LOGIC;�   4   6  <      )           s_axis_tready : out STD_LOGIC;�   3   5  <      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  <      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  <      )           m_axis_tready : in  STD_LOGIC;�   .   0  <      )           m_axis_tlast  : out STD_LOGIC;�   -   /  <      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  <      	    port(�   *   ,  <         component mapper is --{{{�   )   +  <      $   end component slice_2from8; --}}}�   (   *  <      *           rst           : in  STD_LOGIC);�   '   )  <      )           clk           : in  STD_LOGIC;�   %   '  <      )           s_axis_tready : out STD_LOGIC;�   $   &  <      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  <      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  <      )           m_axis_tready : in  STD_LOGIC;�      !  <      )           m_axis_tlast  : out STD_LOGIC;�         <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_2from8 is --{{{�        <      $   end component slice_1from8; --}}}�        <      *           rst           : in  STD_LOGIC);�        <      )           clk           : in  STD_LOGIC;�        <      )           s_axis_tready : out STD_LOGIC;�        <      )           s_axis_tlast  : in  STD_LOGIC;�        <      )           s_axis_tvalid : in  STD_LOGIC;�        <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        <      )           m_axis_tready : in  STD_LOGIC;�        <      )           m_axis_tlast  : out STD_LOGIC;�        <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_1from8 is --{{{�        <      .   signal rst_tb            : STD_LOGIC:= '0';�   
     <      .   signal clk_tb            : STD_LOGIC:= '0';�      
  <      4   signal state   :axiStates := waitingSvalid; --}}}�      	  <      6   type   axiStates is (waitingSvalid, waitingMready);�   w   y          )           s_axis_tready : out STD_LOGIC;�   z   |          0           m_axis_config_tvalid : out STD_LOGIC;�   {   }          0           m_axis_config_tready : in  STD_LOGIC;�   ~   �          *           rst           : in  STD_LOGIC);�   }             )           clk           : in  STD_LOGIC;�   y   {          D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   v   x          )           s_axis_tlast  : in  STD_LOGIC;�   u   w          )           s_axis_tvalid : in  STD_LOGIC;�   t   v          >           s_axis_tdata  : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t          )           m_axis_tready : in  STD_LOGIC;�   q   s          )           m_axis_tlast  : out STD_LOGIC;�   p   r          )           m_axis_tvalid : out STD_LOGIC;�   o   q          =           e_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  	            9        ����                                                                                                                                                                                                                                                                                                                           9   .      9   .       V   .    ^$D     �  9  ;  <      <           rst                  => rst_tb           ); --}}}�  8  :  <      +           clk                  => clk_tb ,�  7  9  <      0           m_axis_config_tready => axis3_tready,�  6  8  <      0           m_axis_config_tvalid => axis3_tvalid,�  5  7  <      /           m_axis_config_tdata  => axis3_tdata,�  4  6  <      1           s_axis_tready        => axis20_tready,�  3  5  <      0           s_axis_tlast         => axis20_tlast,�  2  4  <      1           s_axis_tvalid        => axis20_tvalid,�  1  3  <      0           s_axis_tdata         => axis20_tdata,�  0  2  <      0           m_axis_tready        => axisO_tready,�  /  1  <      /           m_axis_tlast         => axisO_tlast,�  .  0  <      0           m_axis_tvalid        => axisO_tvalid,�  -  /  <      /           m_axis_tdata         => axisO_tdata,�  ,  .  <          port map(  �  *  ,  <      <           rst                  => rst_tb           ); --}}}�  )  +  <      5           clk                  => clk_tb           ,�  (  *  <      1           s_axis_tready        => axis10_tready,�  '  )  <      0           s_axis_tlast         => axis10_tlast,�  &  (  <      1           s_axis_tvalid        => axis10_tvalid,�  %  '  <      0           s_axis_tdata         => axis10_tdata,�  $  &  <      1           m_axis_tready        => axis20_tready,�  #  %  <      0           m_axis_tlast         => axis20_tlast,�  "  $  <      1           m_axis_tvalid        => axis20_tvalid,�  !  #  <      0           m_axis_tdata         => axis20_tdata,�     "  <          port map(  �       <      <           rst                  => rst_tb           ); --}}}�      <      5           clk                  => clk_tb           ,�      <      0           m_axis_config_tready => axis4_tready,�      <      0           m_axis_config_tvalid => axis4_tvalid,�      <      /           m_axis_config_tdata  => axis4_tdata,�      <      2           s_axis_tready        => m1_axis_tready,�      <      1           s_axis_tlast         => m1_axis_tlast,�      <      2           s_axis_tvalid        => m1_axis_tvalid,�      <      1           s_axis_tdata         => m1_axis_tdata,�      <      1           m_axis_tready        => axis10_tready,�      <      0           m_axis_tlast         => axis10_tlast,�      <      1           m_axis_tvalid        => axis10_tvalid,�      <      0           m_axis_tdata         => axis10_tdata,�      <          port map(  �      <      6--           rst           =>rst_tb           ); --}}}�      <      /--           clk           =>clk_tb           ,�      <      *--           s_axis_tready =>axis2_tready,�      <      )--           s_axis_tlast  =>axis2_tlast,�  
    <      *--           s_axis_tvalid =>axis2_tvalid,�  	    <      )--           s_axis_tdata  =>axis2_tdata,�    
  <      *--           m_axis_tready =>axisO_tready,�    	  <      (--           m_axis_tlast  >axisO_tlast,�      <      *--           m_axis_tvalid =>axisO_tvalid,�      <      )--           m_axis_tdata  =>axisO_tdata,�      <      --    port map(  �      <      --             ITER  => 10)�      <      --             N     => 16,�      <      --   generic map(�   �    <      6--           rst           =>rst_tb           ); --}}}�   �     <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m1_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  <      *--           m_axis_tready =>axis2_tready,�   �   �  <      )--           m_axis_tlast  =>axis2_tlast,�   �   �  <      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  <      )--           m_axis_tdata  =>axis2_tdata,�   �   �  <      --    port map(�   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      %   end process axi_master_proc; --}}}�   �   �  <            end if;�   �   �  <               end if;�   �   �  <                  end case;�   �   �  <                        end if;�   �   �  <                           end if;�   �   �  <      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      .                        s1_axis_tready <= '1';�   �   �  <      .                        m1_axis_tvalid <= '0';�   �   �  <                           else�   �   �  <      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  <      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  <      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  <      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  <      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  <      $               when waitingMready =>�   �   �  <                        end if;�   �   �  <      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  <      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  <      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  <      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  <                           end if;�   �   �  <      +                        data2 := data2 + 1;�   �   �  <                           else�   �   �  <      #                        data2 := 0;�   �   �  <      &                     if data2= 15 then�   �   �  <      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  <      )                     bitCounter     := 0;�   �   �  <      *                     s1_axis_tready <='0';�   �   �  <      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  <      $               when waitingSvalid =>�   �   �  <                  case state is�   �   �  <               else�   �   �  <                  data2         := 0;�   �   �  <                  data         := 0;�   �   �  <      .            m1_axis_tdata  <= (others => '0');�   �   �  <      "            m1_axis_tvalid <= '0';�   �   �  <      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  <      "            s1_axis_tready <= '1';�   �   �  <      ,            state          <= waitingSvalid;�   �   �  <               if rst_tb = '0' then�   �   �  <      !      if rising_edge(clk_tb) then�   �   �  <         begin�   �   �  <      ,      variable data2 :natural range 0 to 15;�   �   �  <      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  <      2      variable data :integer range -128 to 127:=0;�   �   �  <      0      variable bitCounter :integer range 0 to 8;�   �   �  <      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  <          rst_tb   <= '1' after 180 ns;�   �   �  <      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  <      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  <      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  <      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  <      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  <      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  <      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  <      )   signal m1_axis_tready: STD_LOGIC:='1';�   �   �  <      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�      �  <      %   end component slice_8from48; --}}}�   ~   �  <      1           rst                  : in  STD_LOGIC);�   }     <      0           clk                  : in  STD_LOGIC;�   {   }  <      0           m_axis_config_tready : in  STD_LOGIC;�   z   |  <      0           m_axis_config_tvalid : out STD_LOGIC;�   y   {  <      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�   w   y  <      0           s_axis_tready        : out STD_LOGIC;�   v   x  <      0           s_axis_tlast         : in  STD_LOGIC;�   u   w  <      0           s_axis_tvalid        : in  STD_LOGIC;�   t   v  <      E           s_axis_tdata         : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  <      0           m_axis_tready        : in  STD_LOGIC;�   q   s  <      0           m_axis_tlast         : out STD_LOGIC;�   p   r  <      0           m_axis_tvalid        : out STD_LOGIC;�   o   q  <      E           e_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);�   n   p  <      	    port(�   m   o  <      #   component slice_8from48 is --{{{�   l   n  <      %   end component join_48from16; --}}}�   k   m  <      *           rst           : in  STD_LOGIC);�   j   l  <      )           clk           : in  STD_LOGIC;�   h   j  <      )           s_axis_tready : out STD_LOGIC;�   g   i  <      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  <      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  <      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  <      )           m_axis_tready : in  STD_LOGIC;�   b   d  <      )           m_axis_tlast  : out STD_LOGIC;�   a   c  <      )           m_axis_tvalid : out STD_LOGIC;�   `   b  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  <      	    port(�   ^   `  <      #   component join_48from16 is --{{{�   ]   _  <      $   end component join_16from8; --}}}�   \   ^  <      *           rst           : in  STD_LOGIC);�   [   ]  <      )           clk           : in  STD_LOGIC;�   Y   [  <      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  <      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  <      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  <      )           s_axis_tready : out STD_LOGIC;�   T   V  <      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  <      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  <      )           m_axis_tready : in  STD_LOGIC;�   O   Q  <      )           m_axis_tlast  : out STD_LOGIC;�   N   P  <      )           m_axis_tvalid : out STD_LOGIC;�   M   O  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  <      	    port(�   K   M  <      "   component join_16from8 is --{{{�   J   L  <         end component cordic; --}}}�   I   K  <      *           rst           : in  STD_LOGIC);�   H   J  <      )           clk           : in  STD_LOGIC;�   F   H  <      )           s_axis_tready : out STD_LOGIC;�   E   G  <      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  <      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  <      )           m_axis_tready : in  STD_LOGIC;�   @   B  <      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  <      )           m_axis_tvalid : out STD_LOGIC;�   >   @  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  <      	    port(�   <   >  <      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  <      9             N     : natural := 16; --Ancho de la palabra�   :   <  <         generic(�   9   ;  <         component cordic is --{{{�   8   :  <         end component mapper; --}}}�   7   9  <      *           rst           : in  STD_LOGIC);�   6   8  <      )           clk           : in  STD_LOGIC;�   4   6  <      )           s_axis_tready : out STD_LOGIC;�   3   5  <      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  <      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  <      )           m_axis_tready : in  STD_LOGIC;�   .   0  <      )           m_axis_tlast  : out STD_LOGIC;�   -   /  <      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  <      	    port(�   *   ,  <         component mapper is --{{{�   )   +  <      $   end component slice_2from8; --}}}�   (   *  <      *           rst           : in  STD_LOGIC);�   '   )  <      )           clk           : in  STD_LOGIC;�   %   '  <      )           s_axis_tready : out STD_LOGIC;�   $   &  <      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  <      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  <      )           m_axis_tready : in  STD_LOGIC;�      !  <      )           m_axis_tlast  : out STD_LOGIC;�         <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_2from8 is --{{{�        <      $   end component slice_1from8; --}}}�        <      *           rst           : in  STD_LOGIC);�        <      )           clk           : in  STD_LOGIC;�        <      )           s_axis_tready : out STD_LOGIC;�        <      )           s_axis_tlast  : in  STD_LOGIC;�        <      )           s_axis_tvalid : in  STD_LOGIC;�        <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        <      )           m_axis_tready : in  STD_LOGIC;�        <      )           m_axis_tlast  : out STD_LOGIC;�        <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_1from8 is --{{{�        <      .   signal rst_tb            : STD_LOGIC:= '0';�   
     <      .   signal clk_tb            : STD_LOGIC:= '0';�      
  <      4   signal state   :axiStates := waitingSvalid; --}}}�      	  <      6   type   axiStates is (waitingSvalid, waitingMready);�  8  :          5           clk                  => clk_tb           ,5�_�                :        ����                                                                                                                                                                                                                                                                                                                           :          :           V        ^$D	     �  9  ;  <      ;           rst                  => rst_tb           );--}}}�  8  :  <      +           clk                  => clk_tb ,�  7  9  <      0           m_axis_config_tready => axis3_tready,�  6  8  <      0           m_axis_config_tvalid => axis3_tvalid,�  5  7  <      /           m_axis_config_tdata  => axis3_tdata,�  4  6  <      1           s_axis_tready        => axis20_tready,�  3  5  <      0           s_axis_tlast         => axis20_tlast,�  2  4  <      1           s_axis_tvalid        => axis20_tvalid,�  1  3  <      0           s_axis_tdata         => axis20_tdata,�  0  2  <      0           m_axis_tready        => axisO_tready,�  /  1  <      /           m_axis_tlast         => axisO_tlast,�  .  0  <      0           m_axis_tvalid        => axisO_tvalid,�  -  /  <      /           m_axis_tdata         => axisO_tdata,�  ,  .  <          port map(  �  *  ,  <      <           rst                  => rst_tb           ); --}}}�  )  +  <      5           clk                  => clk_tb           ,�  (  *  <      1           s_axis_tready        => axis10_tready,�  '  )  <      0           s_axis_tlast         => axis10_tlast,�  &  (  <      1           s_axis_tvalid        => axis10_tvalid,�  %  '  <      0           s_axis_tdata         => axis10_tdata,�  $  &  <      1           m_axis_tready        => axis20_tready,�  #  %  <      0           m_axis_tlast         => axis20_tlast,�  "  $  <      1           m_axis_tvalid        => axis20_tvalid,�  !  #  <      0           m_axis_tdata         => axis20_tdata,�     "  <          port map(  �       <      <           rst                  => rst_tb           ); --}}}�      <      5           clk                  => clk_tb           ,�      <      0           m_axis_config_tready => axis4_tready,�      <      0           m_axis_config_tvalid => axis4_tvalid,�      <      /           m_axis_config_tdata  => axis4_tdata,�      <      2           s_axis_tready        => m1_axis_tready,�      <      1           s_axis_tlast         => m1_axis_tlast,�      <      2           s_axis_tvalid        => m1_axis_tvalid,�      <      1           s_axis_tdata         => m1_axis_tdata,�      <      1           m_axis_tready        => axis10_tready,�      <      0           m_axis_tlast         => axis10_tlast,�      <      1           m_axis_tvalid        => axis10_tvalid,�      <      0           m_axis_tdata         => axis10_tdata,�      <          port map(  �      <      6--           rst           =>rst_tb           ); --}}}�      <      /--           clk           =>clk_tb           ,�      <      *--           s_axis_tready =>axis2_tready,�      <      )--           s_axis_tlast  =>axis2_tlast,�  
    <      *--           s_axis_tvalid =>axis2_tvalid,�  	    <      )--           s_axis_tdata  =>axis2_tdata,�    
  <      *--           m_axis_tready =>axisO_tready,�    	  <      (--           m_axis_tlast  >axisO_tlast,�      <      *--           m_axis_tvalid =>axisO_tvalid,�      <      )--           m_axis_tdata  =>axisO_tdata,�      <      --    port map(  �      <      --             ITER  => 10)�      <      --             N     => 16,�      <      --   generic map(�   �    <      6--           rst           =>rst_tb           ); --}}}�   �     <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m1_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  <      *--           m_axis_tready =>axis2_tready,�   �   �  <      )--           m_axis_tlast  =>axis2_tlast,�   �   �  <      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  <      )--           m_axis_tdata  =>axis2_tdata,�   �   �  <      --    port map(�   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      %   end process axi_master_proc; --}}}�   �   �  <            end if;�   �   �  <               end if;�   �   �  <                  end case;�   �   �  <                        end if;�   �   �  <                           end if;�   �   �  <      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      .                        s1_axis_tready <= '1';�   �   �  <      .                        m1_axis_tvalid <= '0';�   �   �  <                           else�   �   �  <      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  <      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  <      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  <      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  <      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  <      $               when waitingMready =>�   �   �  <                        end if;�   �   �  <      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  <      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  <      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  <      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  <                           end if;�   �   �  <      +                        data2 := data2 + 1;�   �   �  <                           else�   �   �  <      #                        data2 := 0;�   �   �  <      &                     if data2= 15 then�   �   �  <      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  <      )                     bitCounter     := 0;�   �   �  <      *                     s1_axis_tready <='0';�   �   �  <      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  <      $               when waitingSvalid =>�   �   �  <                  case state is�   �   �  <               else�   �   �  <                  data2         := 0;�   �   �  <                  data         := 0;�   �   �  <      .            m1_axis_tdata  <= (others => '0');�   �   �  <      "            m1_axis_tvalid <= '0';�   �   �  <      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  <      "            s1_axis_tready <= '1';�   �   �  <      ,            state          <= waitingSvalid;�   �   �  <               if rst_tb = '0' then�   �   �  <      !      if rising_edge(clk_tb) then�   �   �  <         begin�   �   �  <      ,      variable data2 :natural range 0 to 15;�   �   �  <      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  <      2      variable data :integer range -128 to 127:=0;�   �   �  <      0      variable bitCounter :integer range 0 to 8;�   �   �  <      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  <          rst_tb   <= '1' after 180 ns;�   �   �  <      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  <      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  <      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  <      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  <      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  <      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  <      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  <      )   signal m1_axis_tready: STD_LOGIC:='1';�   �   �  <      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�      �  <      %   end component slice_8from48; --}}}�   ~   �  <      1           rst                  : in  STD_LOGIC);�   }     <      0           clk                  : in  STD_LOGIC;�   {   }  <      0           m_axis_config_tready : in  STD_LOGIC;�   z   |  <      0           m_axis_config_tvalid : out STD_LOGIC;�   y   {  <      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�   w   y  <      0           s_axis_tready        : out STD_LOGIC;�   v   x  <      0           s_axis_tlast         : in  STD_LOGIC;�   u   w  <      0           s_axis_tvalid        : in  STD_LOGIC;�   t   v  <      E           s_axis_tdata         : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  <      0           m_axis_tready        : in  STD_LOGIC;�   q   s  <      0           m_axis_tlast         : out STD_LOGIC;�   p   r  <      0           m_axis_tvalid        : out STD_LOGIC;�   o   q  <      E           e_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);�   n   p  <      	    port(�   m   o  <      #   component slice_8from48 is --{{{�   l   n  <      %   end component join_48from16; --}}}�   k   m  <      *           rst           : in  STD_LOGIC);�   j   l  <      )           clk           : in  STD_LOGIC;�   h   j  <      )           s_axis_tready : out STD_LOGIC;�   g   i  <      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  <      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  <      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  <      )           m_axis_tready : in  STD_LOGIC;�   b   d  <      )           m_axis_tlast  : out STD_LOGIC;�   a   c  <      )           m_axis_tvalid : out STD_LOGIC;�   `   b  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  <      	    port(�   ^   `  <      #   component join_48from16 is --{{{�   ]   _  <      $   end component join_16from8; --}}}�   \   ^  <      *           rst           : in  STD_LOGIC);�   [   ]  <      )           clk           : in  STD_LOGIC;�   Y   [  <      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  <      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  <      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  <      )           s_axis_tready : out STD_LOGIC;�   T   V  <      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  <      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  <      )           m_axis_tready : in  STD_LOGIC;�   O   Q  <      )           m_axis_tlast  : out STD_LOGIC;�   N   P  <      )           m_axis_tvalid : out STD_LOGIC;�   M   O  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  <      	    port(�   K   M  <      "   component join_16from8 is --{{{�   J   L  <         end component cordic; --}}}�   I   K  <      *           rst           : in  STD_LOGIC);�   H   J  <      )           clk           : in  STD_LOGIC;�   F   H  <      )           s_axis_tready : out STD_LOGIC;�   E   G  <      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  <      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  <      )           m_axis_tready : in  STD_LOGIC;�   @   B  <      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  <      )           m_axis_tvalid : out STD_LOGIC;�   >   @  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  <      	    port(�   <   >  <      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  <      9             N     : natural := 16; --Ancho de la palabra�   :   <  <         generic(�   9   ;  <         component cordic is --{{{�   8   :  <         end component mapper; --}}}�   7   9  <      *           rst           : in  STD_LOGIC);�   6   8  <      )           clk           : in  STD_LOGIC;�   4   6  <      )           s_axis_tready : out STD_LOGIC;�   3   5  <      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  <      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  <      )           m_axis_tready : in  STD_LOGIC;�   .   0  <      )           m_axis_tlast  : out STD_LOGIC;�   -   /  <      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  <      	    port(�   *   ,  <         component mapper is --{{{�   )   +  <      $   end component slice_2from8; --}}}�   (   *  <      *           rst           : in  STD_LOGIC);�   '   )  <      )           clk           : in  STD_LOGIC;�   %   '  <      )           s_axis_tready : out STD_LOGIC;�   $   &  <      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  <      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  <      )           m_axis_tready : in  STD_LOGIC;�      !  <      )           m_axis_tlast  : out STD_LOGIC;�         <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_2from8 is --{{{�        <      $   end component slice_1from8; --}}}�        <      *           rst           : in  STD_LOGIC);�        <      )           clk           : in  STD_LOGIC;�        <      )           s_axis_tready : out STD_LOGIC;�        <      )           s_axis_tlast  : in  STD_LOGIC;�        <      )           s_axis_tvalid : in  STD_LOGIC;�        <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        <      )           m_axis_tready : in  STD_LOGIC;�        <      )           m_axis_tlast  : out STD_LOGIC;�        <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_1from8 is --{{{�        <      .   signal rst_tb            : STD_LOGIC:= '0';�   
     <      .   signal clk_tb            : STD_LOGIC:= '0';�      
  <      4   signal state   :axiStates := waitingSvalid; --}}}�      	  <      6   type   axiStates is (waitingSvalid, waitingMready);�  9  ;          <           rst                  => rst_tb           ); --}}}5�_�                :   *    ����                                                                                                                                                                                                                                                                                                                           :          :           V        ^$D     �  9  ;  <      ;           rst                  => rst_tb           );--}}}5�_�                :   ,    ����                                                                                                                                                                                                                                                                                                                           :          :           V        ^$D   � �  9  ;  <      1           rst                  => rst_tb );--}}}5�_�                *        ����                                                                                                                                                                                                                                                                                                                           *         *          V       ^$D     �  9  ;  <      2           rst                  => rst_tb ); --}}}�  8  :  <      +           clk                  => clk_tb ,�  7  9  <      0           m_axis_config_tready => axis3_tready,�  6  8  <      0           m_axis_config_tvalid => axis3_tvalid,�  5  7  <      /           m_axis_config_tdata  => axis3_tdata,�  4  6  <      1           s_axis_tready        => axis20_tready,�  3  5  <      0           s_axis_tlast         => axis20_tlast,�  2  4  <      1           s_axis_tvalid        => axis20_tvalid,�  1  3  <      0           s_axis_tdata         => axis20_tdata,�  0  2  <      0           m_axis_tready        => axisO_tready,�  /  1  <      /           m_axis_tlast         => axisO_tlast,�  .  0  <      0           m_axis_tvalid        => axisO_tvalid,�  -  /  <      /           m_axis_tdata         => axisO_tdata,�  ,  .  <          port map(  �  *  ,  <      <           rst                  => rst_tb           ); --}}}�  )  +  <      +           clk                  => clk_tb ,�  (  *  <      1           s_axis_tready        => axis10_tready,�  '  )  <      0           s_axis_tlast         => axis10_tlast,�  &  (  <      1           s_axis_tvalid        => axis10_tvalid,�  %  '  <      0           s_axis_tdata         => axis10_tdata,�  $  &  <      1           m_axis_tready        => axis20_tready,�  #  %  <      0           m_axis_tlast         => axis20_tlast,�  "  $  <      1           m_axis_tvalid        => axis20_tvalid,�  !  #  <      0           m_axis_tdata         => axis20_tdata,�     "  <          port map(  �       <      <           rst                  => rst_tb           ); --}}}�      <      5           clk                  => clk_tb           ,�      <      0           m_axis_config_tready => axis4_tready,�      <      0           m_axis_config_tvalid => axis4_tvalid,�      <      /           m_axis_config_tdata  => axis4_tdata,�      <      2           s_axis_tready        => m1_axis_tready,�      <      1           s_axis_tlast         => m1_axis_tlast,�      <      2           s_axis_tvalid        => m1_axis_tvalid,�      <      1           s_axis_tdata         => m1_axis_tdata,�      <      1           m_axis_tready        => axis10_tready,�      <      0           m_axis_tlast         => axis10_tlast,�      <      1           m_axis_tvalid        => axis10_tvalid,�      <      0           m_axis_tdata         => axis10_tdata,�      <          port map(  �      <      6--           rst           =>rst_tb           ); --}}}�      <      /--           clk           =>clk_tb           ,�      <      *--           s_axis_tready =>axis2_tready,�      <      )--           s_axis_tlast  =>axis2_tlast,�  
    <      *--           s_axis_tvalid =>axis2_tvalid,�  	    <      )--           s_axis_tdata  =>axis2_tdata,�    
  <      *--           m_axis_tready =>axisO_tready,�    	  <      (--           m_axis_tlast  >axisO_tlast,�      <      *--           m_axis_tvalid =>axisO_tvalid,�      <      )--           m_axis_tdata  =>axisO_tdata,�      <      --    port map(  �      <      --             ITER  => 10)�      <      --             N     => 16,�      <      --   generic map(�   �    <      6--           rst           =>rst_tb           ); --}}}�   �     <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m1_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  <      *--           m_axis_tready =>axis2_tready,�   �   �  <      )--           m_axis_tlast  =>axis2_tlast,�   �   �  <      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  <      )--           m_axis_tdata  =>axis2_tdata,�   �   �  <      --    port map(�   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      6--           rst           =>rst_tb           ); --}}}�   �   �  <      /--           clk           =>clk_tb           ,�   �   �  <      ,--           s_axis_tready =>m3_axis_tready,�   �   �  <      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  <      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  <      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  <      ,--           m_axis_tready =>s3_axis_tready,�   �   �  <      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  <      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  <      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  <      --    port map(  �   �   �  <      %   end process axi_master_proc; --}}}�   �   �  <            end if;�   �   �  <               end if;�   �   �  <                  end case;�   �   �  <                        end if;�   �   �  <                           end if;�   �   �  <      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      .                        s1_axis_tready <= '1';�   �   �  <      .                        m1_axis_tvalid <= '0';�   �   �  <                           else�   �   �  <      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  <      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  <      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  <      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  <      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  <      $               when waitingMready =>�   �   �  <                        end if;�   �   �  <      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  <      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  <      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  <      D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  <      M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  <                           end if;�   �   �  <      +                        data2 := data2 + 1;�   �   �  <                           else�   �   �  <      #                        data2 := 0;�   �   �  <      &                     if data2= 15 then�   �   �  <      E                     data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  <      )                     bitCounter     := 0;�   �   �  <      *                     s1_axis_tready <='0';�   �   �  <      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  <      $               when waitingSvalid =>�   �   �  <                  case state is�   �   �  <               else�   �   �  <                  data2         := 0;�   �   �  <                  data         := 0;�   �   �  <      .            m1_axis_tdata  <= (others => '0');�   �   �  <      "            m1_axis_tvalid <= '0';�   �   �  <      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  <      "            s1_axis_tready <= '1';�   �   �  <      ,            state          <= waitingSvalid;�   �   �  <               if rst_tb = '0' then�   �   �  <      !      if rising_edge(clk_tb) then�   �   �  <         begin�   �   �  <      ,      variable data2 :natural range 0 to 15;�   �   �  <      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  <      2      variable data :integer range -128 to 127:=0;�   �   �  <      0      variable bitCounter :integer range 0 to 8;�   �   �  <      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  <          rst_tb   <= '1' after 180 ns;�   �   �  <      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  <      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  <      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  <      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  <      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  <      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  <      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  <      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  <      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  <      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  <      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  <      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  <      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  <      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  <      )   signal m1_axis_tready: STD_LOGIC:='1';�   �   �  <      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   �   �  <      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   �   �  <      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�      �  <      %   end component slice_8from48; --}}}�   ~   �  <      1           rst                  : in  STD_LOGIC);�   }     <      0           clk                  : in  STD_LOGIC;�   {   }  <      0           m_axis_config_tready : in  STD_LOGIC;�   z   |  <      0           m_axis_config_tvalid : out STD_LOGIC;�   y   {  <      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�   w   y  <      0           s_axis_tready        : out STD_LOGIC;�   v   x  <      0           s_axis_tlast         : in  STD_LOGIC;�   u   w  <      0           s_axis_tvalid        : in  STD_LOGIC;�   t   v  <      E           s_axis_tdata         : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  <      0           m_axis_tready        : in  STD_LOGIC;�   q   s  <      0           m_axis_tlast         : out STD_LOGIC;�   p   r  <      0           m_axis_tvalid        : out STD_LOGIC;�   o   q  <      E           e_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);�   n   p  <      	    port(�   m   o  <      #   component slice_8from48 is --{{{�   l   n  <      %   end component join_48from16; --}}}�   k   m  <      *           rst           : in  STD_LOGIC);�   j   l  <      )           clk           : in  STD_LOGIC;�   h   j  <      )           s_axis_tready : out STD_LOGIC;�   g   i  <      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  <      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  <      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  <      )           m_axis_tready : in  STD_LOGIC;�   b   d  <      )           m_axis_tlast  : out STD_LOGIC;�   a   c  <      )           m_axis_tvalid : out STD_LOGIC;�   `   b  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  <      	    port(�   ^   `  <      #   component join_48from16 is --{{{�   ]   _  <      $   end component join_16from8; --}}}�   \   ^  <      *           rst           : in  STD_LOGIC);�   [   ]  <      )           clk           : in  STD_LOGIC;�   Y   [  <      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  <      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  <      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  <      )           s_axis_tready : out STD_LOGIC;�   T   V  <      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  <      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  <      )           m_axis_tready : in  STD_LOGIC;�   O   Q  <      )           m_axis_tlast  : out STD_LOGIC;�   N   P  <      )           m_axis_tvalid : out STD_LOGIC;�   M   O  <      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  <      	    port(�   K   M  <      "   component join_16from8 is --{{{�   J   L  <         end component cordic; --}}}�   I   K  <      *           rst           : in  STD_LOGIC);�   H   J  <      )           clk           : in  STD_LOGIC;�   F   H  <      )           s_axis_tready : out STD_LOGIC;�   E   G  <      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  <      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  <      )           m_axis_tready : in  STD_LOGIC;�   @   B  <      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  <      )           m_axis_tvalid : out STD_LOGIC;�   >   @  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  <      	    port(�   <   >  <      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  <      9             N     : natural := 16; --Ancho de la palabra�   :   <  <         generic(�   9   ;  <         component cordic is --{{{�   8   :  <         end component mapper; --}}}�   7   9  <      *           rst           : in  STD_LOGIC);�   6   8  <      )           clk           : in  STD_LOGIC;�   4   6  <      )           s_axis_tready : out STD_LOGIC;�   3   5  <      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  <      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  <      )           m_axis_tready : in  STD_LOGIC;�   .   0  <      )           m_axis_tlast  : out STD_LOGIC;�   -   /  <      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  <      	    port(�   *   ,  <         component mapper is --{{{�   )   +  <      $   end component slice_2from8; --}}}�   (   *  <      *           rst           : in  STD_LOGIC);�   '   )  <      )           clk           : in  STD_LOGIC;�   %   '  <      )           s_axis_tready : out STD_LOGIC;�   $   &  <      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  <      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  <      )           m_axis_tready : in  STD_LOGIC;�      !  <      )           m_axis_tlast  : out STD_LOGIC;�         <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_2from8 is --{{{�        <      $   end component slice_1from8; --}}}�        <      *           rst           : in  STD_LOGIC);�        <      )           clk           : in  STD_LOGIC;�        <      )           s_axis_tready : out STD_LOGIC;�        <      )           s_axis_tlast  : in  STD_LOGIC;�        <      )           s_axis_tvalid : in  STD_LOGIC;�        <      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        <      )           m_axis_tready : in  STD_LOGIC;�        <      )           m_axis_tlast  : out STD_LOGIC;�        <      )           m_axis_tvalid : out STD_LOGIC;�        <      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        <      	    port(�        <      "   component slice_1from8 is --{{{�        <      .   signal rst_tb            : STD_LOGIC:= '0';�   
     <      .   signal clk_tb            : STD_LOGIC:= '0';�      
  <      4   signal state   :axiStates := waitingSvalid; --}}}�      	  <      6   type   axiStates is (waitingSvalid, waitingMready);�  )  +          5           clk                  => clk_tb           ,5�_�                 p       ����                                                                                                                                                                                                                                                                                                                           *         *          V       ^$D.   � �   o   q  <      E           e_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);5�_�                 �        ����                                                                                                                                                                                                                                                                                                                           *         *          V       ^$E�     �   �   �           5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F     �   �   �  ;      &                     if data2= 15 then   #                        data2 := 0;                        else   +                        data2 := data2 + 1;                        end if;   M                     --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));   D                     m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  ;      E                     data1 := std_logic_vector(to_unsigned(data2,4));5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F     �   �   �  <                           �   �   �  ;    5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F#     �   �   �  <      O  --                   --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F#     �   �   �  <      N --                   --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F#     �   �   �  <      M--                   --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F#     �   �   �  <      L-                   --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F&     �   �   �  <      K                   --m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F&     �   �   �  <      J                   -m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F'     �   �   �          &                     m1_axis_tdata <= 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^$F*     �   �   �  ;      I                   m1_axis_tdata  <= std_logic_vector(to_signed(data,8));5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$F9     �  8  :  ;      2           rst                  => rst_tb ); --}}}�  7  9  ;      +           clk                  => clk_tb ,�  6  8  ;      0           m_axis_config_tready => axis3_tready,�  5  7  ;      0           m_axis_config_tvalid => axis3_tvalid,�  4  6  ;      /           m_axis_config_tdata  => axis3_tdata,�  3  5  ;      1           s_axis_tready        => axis20_tready,�  2  4  ;      0           s_axis_tlast         => axis20_tlast,�  1  3  ;      1           s_axis_tvalid        => axis20_tvalid,�  0  2  ;      0           s_axis_tdata         => axis20_tdata,�  /  1  ;      0           m_axis_tready        => axisO_tready,�  .  0  ;      /           m_axis_tlast         => axisO_tlast,�  -  /  ;      0           m_axis_tvalid        => axisO_tvalid,�  ,  .  ;      /           m_axis_tdata         => axisO_tdata,�  +  -  ;          port map(  �  )  +  ;      <           rst                  => rst_tb           ); --}}}�  (  *  ;      +           clk                  => clk_tb ,�  '  )  ;      1           s_axis_tready        => axis10_tready,�  &  (  ;      0           s_axis_tlast         => axis10_tlast,�  %  '  ;      1           s_axis_tvalid        => axis10_tvalid,�  $  &  ;      0           s_axis_tdata         => axis10_tdata,�  #  %  ;      1           m_axis_tready        => axis20_tready,�  "  $  ;      0           m_axis_tlast         => axis20_tlast,�  !  #  ;      1           m_axis_tvalid        => axis20_tvalid,�     "  ;      0           m_axis_tdata         => axis20_tdata,�    !  ;          port map(  �      ;      <           rst                  => rst_tb           ); --}}}�      ;      5           clk                  => clk_tb           ,�      ;      0           m_axis_config_tready => axis4_tready,�      ;      0           m_axis_config_tvalid => axis4_tvalid,�      ;      /           m_axis_config_tdata  => axis4_tdata,�      ;      2           s_axis_tready        => m1_axis_tready,�      ;      1           s_axis_tlast         => m1_axis_tlast,�      ;      2           s_axis_tvalid        => m1_axis_tvalid,�      ;      1           s_axis_tdata         => m1_axis_tdata,�      ;      1           m_axis_tready        => axis10_tready,�      ;      0           m_axis_tlast         => axis10_tlast,�      ;      1           m_axis_tvalid        => axis10_tvalid,�      ;      0           m_axis_tdata         => axis10_tdata,�      ;          port map(  �      ;      6--           rst           =>rst_tb           ); --}}}�      ;      /--           clk           =>clk_tb           ,�      ;      *--           s_axis_tready =>axis2_tready,�  
    ;      )--           s_axis_tlast  =>axis2_tlast,�  	    ;      *--           s_axis_tvalid =>axis2_tvalid,�    
  ;      )--           s_axis_tdata  =>axis2_tdata,�    	  ;      *--           m_axis_tready =>axisO_tready,�      ;      (--           m_axis_tlast  >axisO_tlast,�      ;      *--           m_axis_tvalid =>axisO_tvalid,�      ;      )--           m_axis_tdata  =>axisO_tdata,�      ;      --    port map(  �      ;      --             ITER  => 10)�      ;      --             N     => 16,�       ;      --   generic map(�   �     ;      6--           rst           =>rst_tb           ); --}}}�   �   �  ;      /--           clk           =>clk_tb           ,�   �   �  ;      ,--           s_axis_tready =>m1_axis_tready,�   �   �  ;      +--           s_axis_tlast  =>m1_axis_tlast,�   �   �  ;      ,--           s_axis_tvalid =>m1_axis_tvalid,�   �   �  ;      +--           s_axis_tdata  =>m1_axis_tdata,�   �   �  ;      *--           m_axis_tready =>axis2_tready,�   �   �  ;      )--           m_axis_tlast  =>axis2_tlast,�   �   �  ;      *--           m_axis_tvalid =>axis2_tvalid,�   �   �  ;      )--           m_axis_tdata  =>axis2_tdata,�   �   �  ;      --    port map(�   �   �  ;      6--           rst           =>rst_tb           ); --}}}�   �   �  ;      /--           clk           =>clk_tb           ,�   �   �  ;      ,--           s_axis_tready =>m3_axis_tready,�   �   �  ;      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  ;      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  ;      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  ;      ,--           m_axis_tready =>s3_axis_tready,�   �   �  ;      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  ;      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  ;      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  ;      --    port map(  �   �   �  ;      6--           rst           =>rst_tb           ); --}}}�   �   �  ;      /--           clk           =>clk_tb           ,�   �   �  ;      ,--           s_axis_tready =>m3_axis_tready,�   �   �  ;      +--           s_axis_tlast  =>m3_axis_tlast,�   �   �  ;      ,--           s_axis_tvalid =>m3_axis_tvalid,�   �   �  ;      +--           s_axis_tdata  =>m3_axis_tdata,�   �   �  ;      ,--           m_axis_tready =>s3_axis_tready,�   �   �  ;      +--           m_axis_tlast  =>s3_axis_tlast,�   �   �  ;      ,--           m_axis_tvalid =>s3_axis_tvalid,�   �   �  ;      +--           m_axis_tdata  =>s3_axis_tdata,�   �   �  ;      --    port map(  �   �   �  ;      %   end process axi_master_proc; --}}}�   �   �  ;            end if;�   �   �  ;               end if;�   �   �  ;                  end case;�   �   �  ;                        end if;�   �   �  ;                           end if;�   �   �  ;      �                        state          <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   �   �  ;      .                        s1_axis_tready <= '1';�   �   �  ;      .                        m1_axis_tvalid <= '0';�   �   �  ;                           else�   �   �  ;      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));�   �   �  ;      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);�   �   �  ;      f                     if bitCounter < 2 then                             --perfecto, porque bit voy?   �   �   �  ;      Q                     bitCounter := bitCounter+1;                     --incremento�   �   �  ;      q                  if m1_axis_tready= '1' then                           --lo puedo empezar a mandar al otro lado?�   �   �  ;      $               when waitingMready =>�   �   �  ;                        end if;�   �   �  ;      ~                     state          <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   �   �  ;      p                     m1_axis_tvalid <= '1';                         --como puedo mandar, le avoso que tengo dato�   �   �  ;      D                     --m1_axis_tdata  <= "0000" & data1(3 downto 0);�   �   �  ;      F  --                   m1_axis_tdata  <= "000000" & data1(1 downto 0);�   �   �  ;      M                       m1_axis_tdata  <= std_logic_vector(to_signed(data,8));�   �   �  ;        --                   end if;�   �   �  ;      -  --                      data2 := data2 + 1;�   �   �  ;        --                   else�   �   �  ;      %  --                      data2 := 0;�   �   �  ;      (  --                   if data2= 15 then�   �   �  ;      G  --                   data1 := std_logic_vector(to_unsigned(data2,4));�   �   �  ;      )                     bitCounter     := 0;�   �   �  ;      *                     s1_axis_tready <='0';�   �   �  ;      r                  if s1_axis_tvalid= '1' then                           --espero e que este listo para enviar algo�   �   �  ;      $               when waitingSvalid =>�   �   �  ;                  case state is�   �   �  ;               else�   �   �  ;                   data2          := 0;�   �   �  ;                   data           := 0;�   �   �  ;      .            m1_axis_tdata  <= (others => '0');�   �   �  ;      "            m1_axis_tvalid <= '0';�   �   �  ;      R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �  ;      "            s1_axis_tready <= '1';�   �   �  ;      ,            state          <= waitingSvalid;�   �   �  ;               if rst_tb = '0' then�   �   �  ;      !      if rising_edge(clk_tb) then�   �   �  ;         begin�   �   �  ;      ,      variable data2 :natural range 0 to 15;�   �   �  ;      4      variable data1 :std_logic_vector (3 downto 0);�   �   �  ;      2      variable data :integer range -128 to 127:=0;�   �   �  ;      0      variable bitCounter :integer range 0 to 8;�   �   �  ;      ,   axi_master_proc:process (clk_tb) is --{{{�   �   �  ;          rst_tb   <= '1' after 180 ns;�   �   �  ;      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   �   �  ;      .   signal axis20_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      (   signal axis20_tlast:  STD_LOGIC:='0';�   �   �  ;      (   signal axis20_tvalid: STD_LOGIC:='0';�   �   �  ;      M   signal axis20_tdata:  STD_LOGIC_VECTOR (47 downto 0):=(others=>'0'); --{{{�   �   �  ;      .   signal axis11_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      (   signal axis11_tlast:  STD_LOGIC:='0';�   �   �  ;      (   signal axis11_tvalid: STD_LOGIC:='0';�   �   �  ;      M   signal axis11_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  ;      .   signal axis10_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      (   signal axis10_tlast:  STD_LOGIC:='0';�   �   �  ;      (   signal axis10_tvalid: STD_LOGIC:='0';�   �   �  ;      M   signal axis10_tdata:  STD_LOGIC_VECTOR (15 downto 0):=(others=>'0'); --{{{�   �   �  ;      .   signal axisO_tready: STD_LOGIC:='1';  --}}}�   �   �  ;      '   signal axisO_tlast:  STD_LOGIC:='0';�   �   �  ;      '   signal axisO_tvalid: STD_LOGIC:='0';�   �   �  ;      L   signal axisO_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{�   �   �  ;      -   signal axis4_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      '   signal axis4_tlast:  STD_LOGIC:='0';�   �   �  ;      '   signal axis4_tvalid: STD_LOGIC:='0';�   �   �  ;      K   signal axis4_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  ;      -   signal axis3_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      '   signal axis3_tlast:  STD_LOGIC:='0';�   �   �  ;      '   signal axis3_tvalid: STD_LOGIC:='0';�   �   �  ;      K   signal axis3_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  ;      -   signal axis2_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      '   signal axis2_tlast:  STD_LOGIC:='0';�   �   �  ;      '   signal axis2_tvalid: STD_LOGIC:='0';�   �   �  ;      K   signal axis2_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�   �   �  ;      /   signal s1_axis_tready: STD_LOGIC:='0'; --}}}�   �   �  ;      )   signal s1_axis_tlast:  STD_LOGIC:='0';�   �   �  ;      )   signal s1_axis_tvalid: STD_LOGIC:='1';�   �   �  ;      H   signal s1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   �   �  ;      )   signal m1_axis_tready: STD_LOGIC:='1';�   �   �  ;      )   signal m1_axis_tlast:  STD_LOGIC:='0';�   �   �  ;      )   signal m1_axis_tvalid: STD_LOGIC:='0';�   �   �  ;      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{�      �  ;      %   end component slice_8from48; --}}}�   ~   �  ;      1           rst                  : in  STD_LOGIC);�   }     ;      0           clk                  : in  STD_LOGIC;�   {   }  ;      0           m_axis_config_tready : in  STD_LOGIC;�   z   |  ;      0           m_axis_config_tvalid : out STD_LOGIC;�   y   {  ;      E           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7  downto 0);�   w   y  ;      0           s_axis_tready        : out STD_LOGIC;�   v   x  ;      0           s_axis_tlast         : in  STD_LOGIC;�   u   w  ;      0           s_axis_tvalid        : in  STD_LOGIC;�   t   v  ;      E           s_axis_tdata         : in  STD_LOGIC_VECTOR (47 downto 0);�   r   t  ;      0           m_axis_tready        : in  STD_LOGIC;�   q   s  ;      0           m_axis_tlast         : out STD_LOGIC;�   p   r  ;      0           m_axis_tvalid        : out STD_LOGIC;�   o   q  ;      E           m_axis_tdata         : out STD_LOGIC_VECTOR (7  downto 0);�   n   p  ;      	    port(�   m   o  ;      #   component slice_8from48 is --{{{�   l   n  ;      %   end component join_48from16; --}}}�   k   m  ;      *           rst           : in  STD_LOGIC);�   j   l  ;      )           clk           : in  STD_LOGIC;�   h   j  ;      )           s_axis_tready : out STD_LOGIC;�   g   i  ;      )           s_axis_tlast  : in  STD_LOGIC;�   f   h  ;      )           s_axis_tvalid : in  STD_LOGIC;�   e   g  ;      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (15 downto 0);�   c   e  ;      )           m_axis_tready : in  STD_LOGIC;�   b   d  ;      )           m_axis_tlast  : out STD_LOGIC;�   a   c  ;      )           m_axis_tvalid : out STD_LOGIC;�   `   b  ;      >           m_axis_tdata  : out STD_LOGIC_VECTOR (47 downto 0);�   _   a  ;      	    port(�   ^   `  ;      #   component join_48from16 is --{{{�   ]   _  ;      $   end component join_16from8; --}}}�   \   ^  ;      *           rst           : in  STD_LOGIC);�   [   ]  ;      )           clk           : in  STD_LOGIC;�   Y   [  ;      0           m_axis_config_tready : in  STD_LOGIC;�   X   Z  ;      0           m_axis_config_tvalid : out STD_LOGIC;�   W   Y  ;      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   U   W  ;      )           s_axis_tready : out STD_LOGIC;�   T   V  ;      )           s_axis_tlast  : in  STD_LOGIC;�   S   U  ;      )           s_axis_tvalid : in  STD_LOGIC;�   R   T  ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   P   R  ;      )           m_axis_tready : in  STD_LOGIC;�   O   Q  ;      )           m_axis_tlast  : out STD_LOGIC;�   N   P  ;      )           m_axis_tvalid : out STD_LOGIC;�   M   O  ;      >           m_axis_tdata  : out STD_LOGIC_VECTOR (15 downto 0);�   L   N  ;      	    port(�   K   M  ;      "   component join_16from8 is --{{{�   J   L  ;         end component cordic; --}}}�   I   K  ;      *           rst           : in  STD_LOGIC);�   H   J  ;      )           clk           : in  STD_LOGIC;�   F   H  ;      )           s_axis_tready : out STD_LOGIC;�   E   G  ;      )           s_axis_tlast  : in  STD_LOGIC;�   D   F  ;      )           s_axis_tvalid : in  STD_LOGIC;�   C   E  ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   A   C  ;      )           m_axis_tready : in  STD_LOGIC;�   @   B  ;      )           m_axis_tlast  : out STD_LOGIC;�   ?   A  ;      )           m_axis_tvalid : out STD_LOGIC;�   >   @  ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   =   ?  ;      	    port(�   <   >  ;      I             ITER  : natural := 10); -- numero de iteraciones por defecto�   ;   =  ;      9             N     : natural := 16; --Ancho de la palabra�   :   <  ;         generic(�   9   ;  ;         component cordic is --{{{�   8   :  ;         end component mapper; --}}}�   7   9  ;      *           rst           : in  STD_LOGIC);�   6   8  ;      )           clk           : in  STD_LOGIC;�   4   6  ;      )           s_axis_tready : out STD_LOGIC;�   3   5  ;      )           s_axis_tlast  : in  STD_LOGIC;�   2   4  ;      )           s_axis_tvalid : in  STD_LOGIC;�   1   3  ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�   /   1  ;      )           m_axis_tready : in  STD_LOGIC;�   .   0  ;      )           m_axis_tlast  : out STD_LOGIC;�   -   /  ;      )           m_axis_tvalid : out STD_LOGIC;�   ,   .  ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   +   -  ;      	    port(�   *   ,  ;         component mapper is --{{{�   )   +  ;      $   end component slice_2from8; --}}}�   (   *  ;      *           rst           : in  STD_LOGIC);�   '   )  ;      )           clk           : in  STD_LOGIC;�   %   '  ;      )           s_axis_tready : out STD_LOGIC;�   $   &  ;      )           s_axis_tlast  : in  STD_LOGIC;�   #   %  ;      )           s_axis_tvalid : in  STD_LOGIC;�   "   $  ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�       "  ;      )           m_axis_tready : in  STD_LOGIC;�      !  ;      )           m_axis_tlast  : out STD_LOGIC;�         ;      )           m_axis_tvalid : out STD_LOGIC;�        ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        ;      	    port(�        ;      "   component slice_2from8 is --{{{�        ;      $   end component slice_1from8; --}}}�        ;      *           rst           : in  STD_LOGIC);�        ;      )           clk           : in  STD_LOGIC;�        ;      )           s_axis_tready : out STD_LOGIC;�        ;      )           s_axis_tlast  : in  STD_LOGIC;�        ;      )           s_axis_tvalid : in  STD_LOGIC;�        ;      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�        ;      )           m_axis_tready : in  STD_LOGIC;�        ;      )           m_axis_tlast  : out STD_LOGIC;�        ;      )           m_axis_tvalid : out STD_LOGIC;�        ;      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�        ;      	    port(�        ;      "   component slice_1from8 is --{{{�        ;      .   signal rst_tb            : STD_LOGIC:= '0';�   
     ;      .   signal clk_tb            : STD_LOGIC:= '0';�      
  ;      4   signal state   :axiStates := waitingSvalid; --}}}�      	  ;      6   type   axiStates is (waitingSvalid, waitingMready);�   �   �          ,            state          <= waitingSvalid;�   �   �                      data         := 0;�   �   �                      data2         := 0;�   �   �          .            m1_axis_tdata  <= (others => '0');�   �   �          "            m1_axis_tvalid <= '0';�   �   �          R            s1_axis_tvalid <= '1'; --que haga de cuentqa que siempre tiene un dato�   �   �          "            s1_axis_tready <= '1';5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$F=     �   �   �  <                             �   �   �  ;    5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$FL     �   �   �  <      N                      --  m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�    "              �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$FM     �   �   �  <      M                      -  m1_axis_tdata<= std_logic_vector(to_signed(data,8));5�_�     #  !      "   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$F]   � �   �   �  <      G                        m1_axis_tdata  <= "000000" & data1(3 downto 2);5�_�  "  $          #   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$F�   � �   �   �  =                             �   �   �  <    5�_�  #  %          $   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$G�     �   �   �          &                       data := data+1;5�_�  $  &          %   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$G�     �   �   �  >    �   �   �  >    5�_�  %  '          &   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$G�     �   �   �          )                       if data = 120 then   '                          data := -120;                          end if;5�_�  &              '   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$G�   � �   �   �  <    �   �   �  <    5�_�             "  !   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^$FN   � �   �   �  <      I                      --  m1_axis_tdata  <= "000000" & data1(3 downto 2);5�_�  	      
      9        ����                                                                                                                                                                                                                                                                                                                           9   .      9   .       V   .    ^$D     �  8  :  <      5eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  	            
  9        ����                                                                                                                                                                                                                                                                                                                           9   .      9   .       V   .    ^$D      �  8  :  <      5eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �  �  �  �  �  2        ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$Ct     �  1  4  5      W           clk           =>clk_tb           , rst           =>rst_tb           ); --}}}5�_�  �              �  2   -    ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$Cu     �  2  3  4    �  1  2  4      D           m_axis_config_tdata  : out STD_LOGIC_VECTOR (7 downto 0);   0           m_axis_config_tvalid : out STD_LOGIC;   0           m_axis_config_tready : in  STD_LOGIC;5�_�  �          �  �  (        ����                                                                                                                                                                                                                                                                                                                              (         (          (    ^$Cd     �  (  )  5    �  '  )  5      's8lice_8from48_inst:slice_8from48 --{{{5�_�  �          �  �     #    ����                                                                                                                                                                                                                                                                                                                              #         #          #    ^$Bu     �      5      0           m_axis_tdata         => fxis10_tdata,   1           m_axis_tvalid        => fxis10_tvalid,   0           m_axis_tlast         => fxis10_tlast,   1           m_axis_tready        => fxis10_tready,5�_�  �          �  �  %   &    ����                                                                                                                                                                                                                                                                                                                           #          %                   ^$2g     �  $  &  5      '           m_axis_config_tready => '1'.5�_�  �          �  �  #       ����                                                                                                                                                                                                                                                                                                                           #         '   &          %    ^$1q     �  "  '  .                 m_axis_tdata  =>,              m_axis_tvalid =>,              m_axis_tlast  =>,              m_axis_tready =>,�  #  $  .    �  "  )  .      (           m_axis_tdata  =>axis0_tdata,,   (           m_axis_tvalid =>axis0_tdata,,   (           m_axis_tlast  =>axis0_tdata,,   (           m_axis_tready =>axis0_tdata,,   4           s_axis_tdata  =>axis20_tdataaxis20_tdata,   )           s_axis_tvalid =>axis20_tvalid,5�_�  �          �  �  #       ����                                                                                                                                                                                                                                                                                                                           #         &   '          &    ^$1f     �  "  (  .                 m_axis_tdata  =>              m_axis_tvalid =>              m_axis_tlast  =>              m_axis_tready =>              s_axis_tdata  =>,�  #  $  .    �  "  (  .      (           m_axis_tdata  =>axis20_tdata,   (           m_axis_tvalid =>axis20_tvalid   (           m_axis_tlast  =>axis20_tlast,   (           m_axis_tready =>axis20_tready              s_axis_tdata  =>,5�_�  �          �  �   �   
    ����                                                                                                                                                                                                                                                                                                                           #         &                 ^$10     �   �   �  .      A   signal :  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');  --{{{5�_�  �      �  �  �         ����                                                                                                                                                                                                                                                                                                                                       '          '    ^$.�     �      .    �       .      6           s_axis_tdata  =>axis10_tdata,m1_axis_tdata,   7           s_axis_tvalid =>axis10_tvalidm1_axis_tvalid,   6           s_axis_tlast  =>axis10_tlast,m1_axis_tlast,   7           s_axis_tready =>axis10_treadym1_axis_tready,   -           clk           =>clk_tb           ,5�_�  �          �  �         ����                                                                                                                                                                                                                                                                                                                                       '          '    ^$.�     �      .    �       .      6           s_axis_tdata  =>maxis10_tdata,1_axis_tdata,   7           s_axis_tvalid =>maxis10_tvalid1_axis_tvalid,   6           s_axis_tlast  =>maxis10_tlast,1_axis_tlast,   7           s_axis_tready =>maxis10_tready1_axis_tready,   -           clk           =>clk_tb           ,5�_�  �      �  �  �   �        ����                                                                                                                                                                                                                                                                                                                            �                     V        ^�G     �   �   �        &--join_16from8_inst:join_16from8 --{{{5�_�  �      �  �  �   �        ����                                                                                                                                                                                                                                                                                                                            �             4       V        ^�?     �   �   �        '--jjoin_16from8_inst:join_16from8 --{{{5�_�  �      �  �  �   �        ����                                                                                                                                                                                                                                                                                                                            �             4       V        ^�3     �   �   �        '--jjoin_16from8_inst:join_16from8 --{{{5�_�  �          �  �   �        ����                                                                                                                                                                                                                                                                                                                            �             4       V        ^�)   � �   �   �        &--join_16from8_inst:join_16from8 --{{{5�_�  P  R      _  Q   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      C                     m1_axis_tdata  <= "00000" & data1(3 downto 0);5�_�  Q  S          R   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      B                     m1_axis_tdata  <= "0000" & data1(3 downto 0);5�_�  R  T          S   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      A                     m1_axis_tdata  <= "0000 & data1(3 downto 0);5�_�  S  U          T   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      @                     m1_axis_tdata  <= "0000& data1(3 downto 0);5�_�  T  V          U   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      ?                     m1_axis_tdata  <= "0000 data1(3 downto 0);5�_�  U  W          V   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      >                     m1_axis_tdata  <= "0000data1(3 downto 0);5�_�  V  X          W   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      =                     m1_axis_tdata  <= "0000ata1(3 downto 0);5�_�  W  Y          X   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      <                     m1_axis_tdata  <= "0000ta1(3 downto 0);5�_�  X  Z          Y   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      ;                     m1_axis_tdata  <= "0000a1(3 downto 0);5�_�  Y  [          Z   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      :                     m1_axis_tdata  <= "00001(3 downto 0);5�_�  Z  \          [   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      9                     m1_axis_tdata  <= "0000(3 downto 0);5�_�  [  ]          \   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      8                     m1_axis_tdata  <= "00003 downto 0);5�_�  \  ^          ]   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      7                     m1_axis_tdata  <= "0000 downto 0);5�_�  ]              ^   �   ,    ����                                                                                                                                                                                                                                                                                                                            }          }          V       ^\     �   �   �   �      6                     m1_axis_tdata  <= "0000downto 0);5�_�  A  C      H  B   �   '    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^.     �   �   �   �      N                     m1_axis_tdata  <= (others=>'0')l"00" & data1(1 downto 0);5�_�  B  D          C   �   4    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^7     �   �   �   �      M                     m1_axis_tdata  <= (others=>'0')"00" & data1(1 downto 0);5�_�  C  E          D   �   4    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^7     �   �   �   �      L                     m1_axis_tdata  <= (others=>'0')00" & data1(1 downto 0);5�_�  D  F          E   �   4    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^7     �   �   �   �      K                     m1_axis_tdata  <= (others=>'0')0" & data1(1 downto 0);5�_�  E  G          F   �   4    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^7     �   �   �   �      J                     m1_axis_tdata  <= (others=>'0')" & data1(1 downto 0);5�_�  F              G   �   4    ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^8   f �   �   �   �      I                     m1_axis_tdata  <= (others=>'0') & data1(1 downto 0);5�_�  :          <  ;   �       ����                                                                                                                                                                                                                                                                                                                            �   '       �   A       v   A    ^�     �   �   �   �    �      �   �      (                     end if;(3 downto 0)5�_�                    F    ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^�     �   ~   �   �      W                     m1_axis_tdata  <= std_logic_vector(to_signed(data(1 downto 0),8));5�_�  i          k  j   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^U�     �   �   �   �      (           maxis_tdata  =>so_axis_tdata,5�_�  V          X  W   
        ����                                                                                                                                                                                                                                                                                                                            
                      V        ^9<     �   	      �       --{{{�   
      �      4   signal clk_tb            : STD_LOGIC:= '0'; --}}}5�_�  G          I  H   :       ����                                                                                                                                                                                                                                                                                                                                                             ^*�     �   :   ;   �    �   9   :   �      M   signal m1_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):=(others=>'0'); --{{{5�_�  9          ;  :   U       ����                                                                                                                                                                                                                                                                                                                            F           H           V        ^z     �   T   V   �      Q            s1_axis_tvalid<= '0'; --que haga de cuentqa que siempre tiene un dato5�_�  4      5  7  6   E        ����                                                                                                                                                                                                                                                                                                                            E   (       H   (       V   (    ^.     �   D   F   �      L   signal so_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0'); {{{�   G   I   �      0   signal so_axis_tready: STD_LOGIC:='0';  --}}}5�_�  4          6  5   F   )    ����                                                                                                                                                                                                                                                                                                                            H   )       F   )       V   )    ^*     �   E   G   �      /   signal so_axis_tvalid: STD_LOGIC:='1'; --{{{�   G   I   �      0   signal so_axis_tready: STD_LOGIC:='0';  --}}}5�_�  $          &  %   �       ����                                                                                                                                                                                                                                                                                                                            �          �   (       v   (    ^q   * �      �   �                 m_axis_tready =>'1',5�_�          $     W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^�   ' �   V   X   �      b                  if '1' then                           --espero e que este listo para enviar algo5�_�                 W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^�   ( �   V   X   �      i                  if '1' = '1'  then                           --espero e que este listo para enviar algo5�_�                  W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^     �   V   X   �      h                  if 1' = '1'  then                           --espero e que este listo para enviar algo5�_�    !              W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^     �   V   X   �      g                  if 1 = '1'  then                           --espero e que este listo para enviar algo5�_�     "          !   W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^     �   V   X   �      f                  if 1 = 1'  then                           --espero e que este listo para enviar algo5�_�  !  #          "   W       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^   ) �   V   X   �      e                  if 1 = 1  then                           --espero e que este listo para enviar algo5�_�  "              #   P       ����                                                                                                                                                                                                                                                                                                                            W          W   $       v   $    ^      �   O   Q   �      Q            s1_axis_tvalid<= '1'; --que haga de cuentqa que siempre tiene un dato5�_�   �           �   �      '    ����                                                                                                                                                                                                                                                                                                                                                       ^�     �         e    �         e      /   signal rst_tb            : STD_LOGIC: = '0';5�_�   �       �   �   �   '        ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   $   &          I   signal s2_axis_tdata:  STD_LOGIC_VECTOR ( 7 downto 0):= (others=>'0');5�_�   �       �   �   �   '        ����                                                                                                                                                                                                                                                                                                                            %           '           V        ^�     �   $   &          I   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0): = (others=>'0');�   %   '          >   signal s2_axis_tvalid: STD_LOGIC:                     ='0';�   &   (          >   signal s2_axis_tlast:  STD_LOGIC:                     ='0';5�_�   �   �       �   �   )        ����                                                                                                                                                                                                                                                                                                                            %           &           V        ^�     �   (   *          "   signal clk_tb : STD_LOGIC:='0';�   )   +          "   signal rst_tb : STD_LOGIC:='0';�      
   e      4   type axiStates is (waitingSvalid, waitingMready);�   	      e      +   signal state:axiStates := waitingSvalid;�         e         component split_1to8 is�         e      	    port(�         e      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         e      )           m_axis_tvalid : out STD_LOGIC;�         e      )           m_axis_tlast  : out STD_LOGIC;�         e      )           m_axis_tready : in  STD_LOGIC;�         e      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         e      )           s_axis_tvalid : in  STD_LOGIC;�         e      )           s_axis_tlast  : in  STD_LOGIC;�         e      )           s_axis_tready : out STD_LOGIC;�         e      )           clk           : in  STD_LOGIC;�         e      *           rst           : in  STD_LOGIC);�         e         end component split_1to8;�         e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         e      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';�         e      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';�          e      -   signal m1_axis_tready_tb : STD_LOGIC:='1';�      !   e      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�       "   e      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';�   !   #   e      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';�   "   $   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�   $   &   e      H   signal s2_axis_tdata:  STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�   %   '   e      )   signal s2_axis_tvalid: STD_LOGIC:='0';�   &   (   e      )   signal s2_axis_tlast:  STD_LOGIC:='0';�   '   )   e      )   signal s2_axis_tready: STD_LOGIC:='1';�   (   *   e      "   signal clk_tb : STD_LOGIC:='0';�   )   +   e      "   signal rst_tb : STD_LOGIC:='0';�   ,   .   e      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   -   /   e          rst_tb   <= '1' after 180 ns;�   /   1   e      &   axi_master_proc:process (clk_tb) is�   0   2   e      0      variable bitCounter :integer range 0 to 8;�   1   3   e      2      variable data :integer range -128 to 127:=0;�   2   4   e         begin�   3   5   e      !      if rising_edge(clk_tb) then�   4   6   e               if rst_tb = '0' then�   5   7   e      +            state         <= waitingSvalid;�   6   8   e      $            s_axis_tready_tb <= '1';�   7   9   e      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato�   8   :   e      $            m_axis_tvalid_tb <= '0';�   9   ;   e      0            m_axis_tdata_tb  <= (others => '0');�   :   <   e                  data  := 0;�   ;   =   e               else�   <   >   e                  case state is�   =   ?   e      $               when waitingSvalid =>�   >   @   e      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   ?   A   e      -                     s_axis_tready_tb <= '0';�   @   B   e      +                     bitCounter       := 0;�   A   C   e      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   B   D   e      J                     data             :=to_integer(to_signed(data + 1,8));�   C   E   e      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   D   F   e      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   E   G   e                        end if;�   F   H   e      $               when waitingMready =>�   G   I   e      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   H   J   e      Q                     bitCounter := bitCounter+1;                     --incremento�   I   K   e      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   J   L   e      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));�   K   M   e      R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   L   N   e                           else�   M   O   e      0                        m_axis_tvalid_tb <= '0';�   N   P   e      0                        s_axis_tready_tb <= '1';�   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   P   R   e                           end if;�   Q   S   e                        end if;�   R   T   e                  end case;�   S   U   e               end if;�   T   V   e            end if;�   U   W   e         end process axi_master_proc;�   X   Z   e          port map(  �   Y   [   e      )           m_axis_tdata  =>s2_axis_tdata,�   Z   \   e      *           m_axis_tvalid =>s2_axis_tvalid,�   [   ]   e      )           m_axis_tlast  =>s2_axis_tlast,�   \   ^   e      *           m_axis_tready =>s2_axis_tready,�   ]   _   e      )           s_axis_tdata  =>m1_axis_tdata,�   ^   `   e      *           s_axis_tvalid =>m1_axis_tvalid,�   _   a   e      )           s_axis_tlast  =>m1_axis_tlast,�   `   b   e      *           s_axis_tready =>m1_axis_tready,�   a   c   e      -           clk           =>clk_tb           ,�   b   d   e      .           rst           =>rst_tb           );5�_�   �       �       �   %        ����                                                                                                                                                                                                                                                                                                                            %           *           V        ^�     �   $   +   e      Heeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   )eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   "eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   "eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�   �           �   �   %        ����                                                                                                                                                                                                                                                                                                                            *           %           V        ^�     �   '   )          J   signal s2_axis_tready: STD_LOGIC:='1'                                 ;�   (   *          J   signal clk_tb : STD_LOGIC:='0'                                        ;�   $   &          J   signal s2_axis_tdata:  STD_LOGIC_VECTOR ( 7 downto 0 ):= (others=>'0');�   %   '          J   signal s2_axis_tvalid: STD_LOGIC:='0'                                 ;�   &   (          J   signal s2_axis_tlast:  STD_LOGIC:='0'                                 ;�   )   +          J   signal rst_tb : STD_LOGIC:='0'                                        ;�      
   e      4   type axiStates is (waitingSvalid, waitingMready);�   	      e      +   signal state:axiStates := waitingSvalid;�         e         component split_1to8 is�         e      	    port(�         e      =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�         e      )           m_axis_tvalid : out STD_LOGIC;�         e      )           m_axis_tlast  : out STD_LOGIC;�         e      )           m_axis_tready : in  STD_LOGIC;�         e      =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         e      )           s_axis_tvalid : in  STD_LOGIC;�         e      )           s_axis_tlast  : in  STD_LOGIC;�         e      )           s_axis_tready : out STD_LOGIC;�         e      )           clk           : in  STD_LOGIC;�         e      *           rst           : in  STD_LOGIC);�         e         end component split_1to8;�         e      K   signal m1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):=(others=>'0');�         e      -   signal m1_axis_tvalid_tb : STD_LOGIC:='0';�         e      -   signal m1_axis_tlast_tb  : STD_LOGIC:='0';�          e      -   signal m1_axis_tready_tb : STD_LOGIC:='1';�      !   e      L   signal s1_axis_tdata_tb  : STD_LOGIC_VECTOR (7 downto 0):= (others=>'0');�       "   e      -   signal s1_axis_tvalid_tb : STD_LOGIC:='1';�   !   #   e      -   signal s1_axis_tlast_tb  : STD_LOGIC:='0';�   "   $   e      -   signal s1_axis_tready_tb : STD_LOGIC:='0';�   $   &   e      J   signal s2_axis_tdata:  STD_LOGIC_VECTOR ( 7 downto 0 ):= (others=>'0');�   %   '   e      J   signal s2_axis_tvalid: STD_LOGIC:='0'                                 ;�   &   (   e      J   signal s2_axis_tlast:  STD_LOGIC:='0'                                 ;�   '   )   e      J   signal s2_axis_tready: STD_LOGIC:='1'                                 ;�   (   *   e      J   signal clk_tb : STD_LOGIC:='0'                                        ;�   )   +   e      J   signal rst_tb : STD_LOGIC:='0'                                        ;�   ,   .   e      /   clk_tb   <= not clk_tb after 100 ns; --10Mhz�   -   /   e          rst_tb   <= '1' after 180 ns;�   /   1   e      &   axi_master_proc:process (clk_tb) is�   0   2   e      0      variable bitCounter :integer range 0 to 8;�   1   3   e      2      variable data :integer range -128 to 127:=0;�   2   4   e         begin�   3   5   e      !      if rising_edge(clk_tb) then�   4   6   e               if rst_tb = '0' then�   5   7   e      +            state         <= waitingSvalid;�   6   8   e      $            s_axis_tready_tb <= '1';�   7   9   e      T            s_axis_tvalid_tb <= '1'; --que haga de cuentqa que siempre tiene un dato�   8   :   e      $            m_axis_tvalid_tb <= '0';�   9   ;   e      0            m_axis_tdata_tb  <= (others => '0');�   :   <   e                  data  := 0;�   ;   =   e               else�   <   >   e                  case state is�   =   ?   e      $               when waitingSvalid =>�   >   @   e      u                  if s_axis_tvalid_tb = '1' then                           --espero e que este listo para enviar algo�   ?   A   e      -                     s_axis_tready_tb <= '0';�   @   B   e      +                     bitCounter       := 0;�   A   C   e      M                     m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   B   D   e      J                     data             :=to_integer(to_signed(data + 1,8));�   C   E   e      r                     m_axis_tvalid_tb <= '1';                         --como puedo mandar, le avoso que tengo dato�   D   F   e      �                     state            <= waitingMready;               --cambio de estado, y le doy un clk para que ponga el dato�   E   G   e                        end if;�   F   H   e      $               when waitingMready =>�   G   I   e      t                  if m_axis_tready_tb = '1' then                           --lo puedo empezar a mandar al otro lado?�   H   J   e      Q                     bitCounter := bitCounter+1;                     --incremento�   I   K   e      f                     if bitCounter < 1 then                             --perfecto, porque bit voy?   �   J   L   e      Z                     m_axis_tdata_tb  <= "10101111";--std_logic_vector(to_signed(data,8));�   K   M   e      R                     --   m_axis_tdata_tb  <= std_logic_vector(to_signed(data,8));�   L   N   e                           else�   M   O   e      0                        m_axis_tvalid_tb <= '0';�   N   P   e      0                        s_axis_tready_tb <= '1';�   O   Q   e      �                        state            <= waitingSvalid;                    --cambio de estado, y le doy un clk para que ponga el dato�   P   R   e                           end if;�   Q   S   e                        end if;�   R   T   e                  end case;�   S   U   e               end if;�   T   V   e            end if;�   U   W   e         end process axi_master_proc;�   X   Z   e          port map(  �   Y   [   e      )           m_axis_tdata  =>s2_axis_tdata,�   Z   \   e      *           m_axis_tvalid =>s2_axis_tvalid,�   [   ]   e      )           m_axis_tlast  =>s2_axis_tlast,�   \   ^   e      *           m_axis_tready =>s2_axis_tready,�   ]   _   e      )           s_axis_tdata  =>m1_axis_tdata,�   ^   `   e      *           s_axis_tvalid =>m1_axis_tvalid,�   _   a   e      )           s_axis_tlast  =>m1_axis_tlast,�   `   b   e      *           s_axis_tready =>m1_axis_tready,�   a   c   e      -           clk           =>clk_tb           ,�   b   d   e      .           rst           =>rst_tb           );5�_�   �           �   �   `   (    ����                                                                                                                                                                                                                                                                                                                            ]          Z                 ^n     �   _   b        5�_�   ~           �      3       ����                                                                                                                                                                                                                                                                                                                            C   )       C   5       v   5    ^    �   2   4   f            variable data :signed:=0;5�_�   U           W   V   G   G    ����                                                                                                                                                                                                                                                                                                                            G   L       G   V       v   V    ^'     �   F   H   `      e                        m_axis_tdata_tb  <= std_logic_vector(to_signed(m_axis_tdata_tb,data'length));5�_�   G           I   H   0       ����                                                                                                                                                                                                                                                                                                                                                             ^P     �   /   1   `      !      if rising_edge(clk)_tb then5�_�                    8       ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^&     �   7   9   e      +            state         <= waitingMready;5�_�                    K   #    ����                                                                                                                                                                                                                                                                                                                            B   7       C   7          7    ^��     �   J   L   e      Z                        m_axis_tdat_tba(0) <= s_axis_tdata(bitCounter);    --pongo el dato5��