Vim�UnDo� aݹ9�~뵼k�i����hP��'��{���o      "architecture Behavioral of 8to1 is                             ^    _�                            ����                                                                                                                                                                                                                                                                                                                                                       ^[     �               #           m_valid : out STD_LOGIC;   #           m_last  : out STD_LOGIC;   #           m_ready : in  STD_LOGIC;       8           s_data  : in  STD_LOGIC_VECTOR (7  downto 0);   #           s_valid : in  STD_LOGIC;   #           s_last  : in  STD_LOGIC;   #           s_ready : out STD_LOGIC;�               8           m_data  : out STD_LOGIC_VECTOR (7  downto 0);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^e     �               (           m_axis_valid : out STD_LOGIC;   (           m_axis_last  : out STD_LOGIC;   (           m_axis_ready : in  STD_LOGIC;       =           s_axis_data  : in  STD_LOGIC_VECTOR (7  downto 0);   (           s_axis_valid : in  STD_LOGIC;   (           s_axis_last  : in  STD_LOGIC;   (           s_axis_ready : out STD_LOGIC;�               =           m_axis_data  : out STD_LOGIC_VECTOR (7  downto 0);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^h     �            	   >           m_axis_udata  : out STD_LOGIC_VECTOR (7  downto 0);   )           m_axis_uvalid : out STD_LOGIC;   )           m_axis_ulast  : out STD_LOGIC;   )           m_axis_uready : in  STD_LOGIC;       >           s_axis_udata  : in  STD_LOGIC_VECTOR (7  downto 0);   )           s_axis_uvalid : in  STD_LOGIC;   )           s_axis_ulast  : in  STD_LOGIC;   )           s_axis_uready : out STD_LOGIC;5�_�                          ����                                                                                                                                                                                                                                                                                                                                                       ^q     �            	   >           m_axis_ydata  : out STD_LOGIC_VECTOR (7  downto 0);   )           m_axis_yvalid : out STD_LOGIC;   )           m_axis_ylast  : out STD_LOGIC;   )           m_axis_yready : in  STD_LOGIC;       >           s_axis_ydata  : in  STD_LOGIC_VECTOR (7  downto 0);   )           s_axis_yvalid : in  STD_LOGIC;   )           s_axis_ylast  : in  STD_LOGIC;   )           s_axis_yready : out STD_LOGIC;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^}    �            	   >           m_axis_edata  : out STD_LOGIC_VECTOR (7  downto 0);   )           m_axis_evalid : out STD_LOGIC;   )           m_axis_elast  : out STD_LOGIC;   )           m_axis_eready : in  STD_LOGIC;       >           s_axis_edata  : in  STD_LOGIC_VECTOR (7  downto 0);   )           s_axis_evalid : in  STD_LOGIC;   )           s_axis_elast  : in  STD_LOGIC;   )           s_axis_eready : out STD_LOGIC;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               entity 8to1 is5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               entity byte2bit8to1 is5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               entity byte2bitto1 is5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               entity byte2bito1 is5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               entity byte2bit1 is5�_�                          ����                                                                                                                                                                                                                                                                                                                                                v       ^�     �               entity byte2bit is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       ^     �               entity byte2bit is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       ^     �               	end 8to1;�             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                v       ^    �               "architecture Behavioral of 8to1 is�             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^�     �               
entity  is5�_�                           ����                                                                                                                                                                                                                                                                                                                                                       ^l     �            	   >           m_axis_edata  : out STD_LOGIC_VECTOR (7  downto 0);   )           m_axis_evalid : out STD_LOGIC;   )           m_axis_elast  : out STD_LOGIC;   )           m_axis_eready : in  STD_LOGIC;       >           s_axis_edata  : in  STD_LOGIC_VECTOR (7  downto 0);   )           s_axis_evalid : in  STD_LOGIC;   )           s_axis_elast  : in  STD_LOGIC;   )           s_axis_eready : out STD_LOGIC;5��