Vim�UnDo� �c�ȈO�jCp���Z2���\-&Z?M�F�   �   0                        if bitCounter = '1' then   �   (  �  �      �  �  �    ^*  � _�      �          �   k   L    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U   � �   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   k   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U)     �   j   l   �      _                                wirez(0) <= std_logic_vector(to_signed(-1800,wirez(0)'length));5�_�  �  �          �   k   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U*     �   j   l   �      ^                                wirez(0) <= std_logic_vector(to_signed(1800,wirez(0)'length));5�_�  �  �          �   k   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U+     �   j   l   �      ]                                wirez(0) <= std_logic_vector(to_signed(800,wirez(0)'length));5�_�  �  �          �   k   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U+     �   j   l   �      \                                wirez(0) <= std_logic_vector(to_signed(00,wirez(0)'length));5�_�  �  �          �   m   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U,   � �   l   n   �      [                                wirez(0) <= std_logic_vector(to_signed(0,wirez(0)'length));5�_�  �  �          �   m   K    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U�   � �   l   n   �      _                                wirez(0) <= std_logic_vector(to_signed(-1800,wirez(0)'length));5�_�  �  �          �   k   G    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U�     �   j   l   �      [                                wirez(0) <= std_logic_vector(to_signed(0,wirez(0)'length));5�_�  �  �          �   k   L    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U�     �   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(180000,wirez(0)'length));5�_�  �  �          �   �   8    ����                                                                                                                                                    Y                                                                                                                                                                      h           h   i       V   (    ^U�   � �   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  �  �          �   d        ����                                                                                                                                                    Y                                                                                                                                                                      d          f          V       ^V�     �   c   d          E                          --wirey(0)(15)          <= s_axis_tdata(7);   N                          --wirey(0)(14 downto 7) <= s_axis_tdata(7 downto 0);   E                          --wirey(0)(6  downto 0) <= (others => '0');5�_�  �  �          �   W        ����                                                                                                                                                    Y                                                                                                                                                                      W          Z          V       ^V�   � �   V   W          9                          --wirex(0)(15)          <= '0';   9                          --wirex(0)(14)          <= '0';   N                          --wirex(0)(13 downto 7) <= s_axis_tdata(6 downto 0);   E                          --wirex(0)(6  downto 0) <= (others => '0');5�_�  �  �          �   u       ����                                                                                                                                                                                                                                                                                                                                                            ^W�   � �   t   v   �      o                  if dv(ITER-1) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                      +          V       ^m�     �      1   �    �          �    �                #             clk   : in  std_logic;   #             rst   : in  std_logic;   #             en_i  : in  std_logic;   #             inv_i : in  std_logic;   9             xi    : in  std_logic_vector (N-1 downto 0);   9             yi    : in  std_logic_vector (N-1 downto 0);   9             zi    : in  std_logic_vector (N-1 downto 0);   9             ci    : in  std_logic_vector (N-1 downto 0);   #             dv_o  : out std_logic;   #             inv_o : out std_logic;   9             xip1  : out std_logic_vector (N-1 downto 0);   9             yip1  : out std_logic_vector (N-1 downto 0);   8             zip1  : out std_logic_vector (N-1 downto 0)5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                       0   (       V       ^m�     �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                                       0   (       V       ^m�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^m�     �   �   �   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);   8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);   "          m_valid : out STD_LOGIC;   "          m_inv   : out STD_LOGIC;   "          m_ready : in  STD_LOGIC;       8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);   8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);   8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);   8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);   "          s_valid : in  STD_LOGIC;   "          s_ready : out STD_LOGIC;   "          s_inv   : in  STD_LOGIC;   "          s_atan  : in  STD_LOGIC;       (          clk           : in  STD_LOGIC;   )          rst           : in  STD_LOGIC);�   �   �   �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �  �      �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   ,       ���    ^m�     �   �   �   �      ;          m_dataX => : out STD_LOGIC_VECTOR (N-1 downto 0);   ;          m_dataY => : out STD_LOGIC_VECTOR (N-1 downto 0);   ;          m_dataZ => : out STD_LOGIC_VECTOR (N-1 downto 0);   %          m_valid => : out STD_LOGIC;   %          m_inv   => : out STD_LOGIC;   %          m_ready => : in  STD_LOGIC;       ;          s_dataX => : in  STD_LOGIC_VECTOR (N-1 downto 0);   ;          s_dataY => : in  STD_LOGIC_VECTOR (N-1 downto 0);   ;          s_dataZ => : in  STD_LOGIC_VECTOR (N-1 downto 0);   ;          s_dataT => : in  STD_LOGIC_VECTOR (N-1 downto 0);   %          s_valid => : in  STD_LOGIC;   %          s_ready => : out STD_LOGIC;   %          s_inv   => : in  STD_LOGIC;   %          s_atan  => : in  STD_LOGIC;       +          clk     =>       : in  STD_LOGIC;   ,          rst     =>       : in  STD_LOGIC);5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   ,       ���    ^m�     �   �   �   �                clk     => 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   ,       ���    ^m�     �   �   �   �                rst     => 5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^m�     �   �   �                           clk   => clk,                    rst   => rst,5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n     �   �   �          *                 en_i  => en      ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n     �   �   �   �                s_ready => 5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n!     �   �   �          *                 en_i  => en      ( j   ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n)     �   �   �          *                 inv_i => inv     ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n*     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n.     �   �   �   �                s_inv   =>    *                 inv_i => inv     ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^n0     �   �   �   �      .          s_inv   => inv_i => inv     ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^n1     �   �   �   �      &          s_inv   =>  inv     ( j   ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n5     �   �   �          *                 xi    => wirex   ( j   ),   *                 yi    => wirey   ( j   ),   *                 zi    => wirez   ( j   ),   *                 ci    => wireLUT ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n8     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   *       ���    ^n>     �   �   �   �                s_dataX =>              s_dataY =>              s_dataZ =>              s_dataT =>    *                 xi    => wirex   ( j   ),�   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n@     �   �   �          *                 xi    => wirex   ( j   ),   *                 yi    => wirey   ( j   ),   *                 zi    => wirez   ( j   ),   *                 ci    => wireLUT ( j   ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^nE     �   �   �          *                 dv_o  => dv      ( j   ),   *                 inv_o => inv     ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^nH     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   *       ���    ^nQ     �   �   �   �                m_valid =>              m_inv   =>              m_ready => �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^nT     �   �   �          *                 dv_o  => dv      ( j   ),   *                 inv_o => inv     ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^nW     �   �   �          *                 xip1  => wirex   ( j+1 ),   *                 yip1  => wirey   ( j+1 ),   )                 zip1  => wirez   ( j+1 )5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^nZ     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �   )          )    ^n`     �   �   �   �                m_dataX =>              m_dataY =>              m_dataZ =>    *                 xip1  => wirex   ( j+1 ),�   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^na     �   �   �          *                 xip1  => wirex   ( j+1 ),   *                 yip1  => wirey   ( j+1 ),   )                 zip1  => wirez   ( j+1 )5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   	       �   	       V   	    ^nl     �   �   �   �         end generate;�   �   �   �               en(j+1)<=dv(j);�   �   �   �                    );�   �   �   �                rst     => rst,�   �   �   �                clk     => clk,�   �   �   �                s_atan  =>�   �   �   �      %          s_inv   => inv     ( j   ),�   �   �   �                s_ready => en(j),�   �   �   �                s_valid =>�   �   �   �      %          s_dataT => wireLUT ( j   ),�   �   �   �      %          s_dataZ => wirez   ( j   ),�   �   �   �      %          s_dataY => wirey   ( j   ),�   �   �   �      %          s_dataX => wirex   ( j   ),�   �   �   �                m_ready =>�   �   �   �      %          m_inv   => inv     ( j+1 ),�   �   �   �      %          m_valid => dv      ( j   ),�   �   �   �      $          m_dataZ => wirez   ( j+1 )�   �   �   �      %          m_dataY => wirey   ( j+1 ),�   �   �   �      %          m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      !                  en ( 0 )<= '0';�   w   y   �      $               when waitingCordic =>�   v   x   �                        end if;�   u   w   �      2                     bitCounter := bitCounter + 1;�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      @                          state                <= waitingCordic;�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   n   p   �      !                          end if;�   m   o   �      :                                wirez(0) <= (others=>'0');�   l   n   �                                else �   k   m   �      $                             end if;�   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   i   k   �      "                             else �   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   g   i   �      8                             if s_axis_tdata(7)='1' then�   f   h   �      ,                          if inv(0)='1' then�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   d   f   �      4                          wirey(0) <= (others=>'0');�   c   e   �      !                        when 1 =>�   b   d   �      !                          end if;�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   [   ]   �      4                          wirex(0) <= (others=>'0');�   Z   \   �      !                        when 0 =>�   Y   [   �      '                     case bitCounter is�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case state is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                    clk     => clk,�   �   �                    s_atan  => �   �   �          %          s_inv   => inv     ( j   ),�   �   �                    s_ready => en(j),�   �   �                    s_valid => �   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),�   �   �                    rst     => rst,�   �   �                    m_ready => �   �   �          %          m_inv   =>inv     ( j+1 ), �   �   �          %          m_valid =>dv      ( j   ), �   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   	       �   	       V   	    ^nm     �   �   �           5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^nq     �   �   �   �         end generate;�   �   �   �               en(j+1)<=dv(j);�   �   �   �                    );�   �   �   �                rst     => rst,�   �   �   �                clk     => clk,�   �   �   �                s_atan  =>�   �   �   �      %          s_inv   => inv     ( j   ),�   �   �   �                s_ready => en(j),�   �   �   �                s_valid =>�   �   �   �      %          s_dataT => wireLUT ( j   ),�   �   �   �      %          s_dataZ => wirez   ( j   ),�   �   �   �      %          s_dataY => wirey   ( j   ),�   �   �   �      %          s_dataX => wirex   ( j   ),�   �   �   �                m_ready =>�   �   �   �      %          m_inv   => inv     ( j+1 ),�   �   �   �      %          m_valid => dv      ( j   ),�   �   �   �      $          m_dataZ => wirez   ( j+1 )�   �   �   �      %          m_dataY => wirey   ( j+1 ),�   �   �   �      %          m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      !                  en ( 0 )<= '0';�   w   y   �      $               when waitingCordic =>�   v   x   �                        end if;�   u   w   �      2                     bitCounter := bitCounter + 1;�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      @                          state                <= waitingCordic;�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   n   p   �      !                          end if;�   m   o   �      :                                wirez(0) <= (others=>'0');�   l   n   �                                else �   k   m   �      $                             end if;�   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   i   k   �      "                             else �   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   g   i   �      8                             if s_axis_tdata(7)='1' then�   f   h   �      ,                          if inv(0)='1' then�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   d   f   �      4                          wirey(0) <= (others=>'0');�   c   e   �      !                        when 1 =>�   b   d   �      !                          end if;�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   [   ]   �      4                          wirex(0) <= (others=>'0');�   Z   \   �      !                        when 0 =>�   Y   [   �      '                     case bitCounter is�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case state is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                    rst     => rst,�   �   �                    clk     => clk,�   �   �                    s_atan  =>�   �   �          %          s_inv   => inv     ( j   ),�   �   �                    s_ready => en(j),�   �   �                    s_valid =>�   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),�   �   �                    m_ready =>�   �   �          %          m_inv   => inv     ( j+1 ),�   �   �          %          m_valid => dv      ( j   ),�   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),�   �   �          %          m_dataX => wirex   ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^ns     �   �   �   �         end generate;�   �   �   �               en(j+1)<=dv(j);�   �   �   �                    );�   �   �   �                rst     => rst,�   �   �   �                clk     => clk,�   �   �   �                s_atan  =>�   �   �   �      %          s_inv   => inv     ( j   ),�   �   �   �      %          s_ready => en      ( j   ),�   �   �   �                s_valid =>�   �   �   �      %          s_dataT => wireLUT ( j   ),�   �   �   �      %          s_dataZ => wirez   ( j   ),�   �   �   �      %          s_dataY => wirey   ( j   ),�   �   �   �      %          s_dataX => wirex   ( j   ),�   �   �   �                m_ready =>�   �   �   �      %          m_inv   => inv     ( j+1 ),�   �   �   �      %          m_valid => dv      ( j   ),�   �   �   �      $          m_dataZ => wirez   ( j+1 )�   �   �   �      %          m_dataY => wirey   ( j+1 ),�   �   �   �      %          m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      !                  en ( 0 )<= '0';�   w   y   �      $               when waitingCordic =>�   v   x   �                        end if;�   u   w   �      2                     bitCounter := bitCounter + 1;�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      @                          state                <= waitingCordic;�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   n   p   �      !                          end if;�   m   o   �      :                                wirez(0) <= (others=>'0');�   l   n   �                                else �   k   m   �      $                             end if;�   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   i   k   �      "                             else �   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   g   i   �      8                             if s_axis_tdata(7)='1' then�   f   h   �      ,                          if inv(0)='1' then�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   d   f   �      4                          wirey(0) <= (others=>'0');�   c   e   �      !                        when 1 =>�   b   d   �      !                          end if;�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   [   ]   �      4                          wirex(0) <= (others=>'0');�   Z   \   �      !                        when 0 =>�   Y   [   �      '                     case bitCounter is�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case state is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          m_valid => dv      ( j   ),�   �   �          %          m_inv   => inv     ( j+1 ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),�   �   �          "          s_ready => en      ( j),�   �   �          %          m_dataX => wirex   ( j+1 ),�   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_inv   => inv     ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          m_valid => dv      ( j   ),�   �   �          %          m_inv   => inv     ( j+1 ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),�   �   �                    s_ready => en(j),�   �   �          %          m_dataX => wirex   ( j+1 ),�   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_inv   => inv     ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^nu     �   �   �   �         end generate;�   �   �   �               en(j+1)<=dv(j);�   �   �   �                    );�   �   �   �                rst     => rst,�   �   �   �                clk     => clk,�   �   �   �                s_atan  =>�   �   �   �      %          s_inv   => inv     ( j   ),�   �   �   �      %          s_ready => en      ( j   ),�   �   �   �                s_valid =>�   �   �   �      %          s_dataT => wireLUT ( j   ),�   �   �   �      %          s_dataZ => wirez   ( j   ),�   �   �   �      %          s_dataY => wirey   ( j   ),�   �   �   �      %          s_dataX => wirex   ( j   ),�   �   �   �                m_ready =>�   �   �   �      %          m_inv   => inv     ( j+1 ),�   �   �   �      %          m_valid => dv      ( j   ),�   �   �   �      $          m_dataZ => wirez   ( j+1 )�   �   �   �      %          m_dataY => wirey   ( j+1 ),�   �   �   �      %          m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      !                  en ( 0 )<= '0';�   w   y   �      $               when waitingCordic =>�   v   x   �                        end if;�   u   w   �      2                     bitCounter := bitCounter + 1;�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      @                          state                <= waitingCordic;�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   n   p   �      !                          end if;�   m   o   �      :                                wirez(0) <= (others=>'0');�   l   n   �                                else �   k   m   �      $                             end if;�   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   i   k   �      "                             else �   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   g   i   �      8                             if s_axis_tdata(7)='1' then�   f   h   �      ,                          if inv(0)='1' then�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   d   f   �      4                          wirey(0) <= (others=>'0');�   c   e   �      !                        when 1 =>�   b   d   �      !                          end if;�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   [   ]   �      4                          wirex(0) <= (others=>'0');�   Z   \   �      !                        when 0 =>�   Y   [   �      '                     case bitCounter is�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case state is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                    rst     => rst,�   �   �                    clk     => clk,�   �   �                    s_atan  =>�   �   �          %          s_inv   => inv     ( j   ),�   �   �          %          s_ready => en      ( j   ),�   �   �                    s_valid =>�   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),�   �   �                    m_ready =>�   �   �          %          m_inv   => inv     ( j+1 ),�   �   �          %          m_valid => dv      ( j   ),�   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),�   �   �          %          m_dataX => wirex   ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^n�     �   �   �           5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �   
       �   
       V   
    ^n�     �   �   �                        );5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n�     �   �   �          	       );�   �   �                    rst     => rst,�   �   �                    clk     => clk,�   �   �                    s_atan  =>�   �   �          %          s_inv   => inv     ( j   ),�   �   �          %          s_ready => en      ( j   ),�   �   �                    s_valid =>�   �   �          %          s_dataT => wireLUT ( j   ),�   �   �          %          s_dataZ => wirez   ( j   ),�   �   �          %          s_dataY => wirey   ( j   ),�   �   �          %          s_dataX => wirex   ( j   ),�   �   �                    m_ready =>�   �   �          %          m_inv   => inv     ( j+1 ),�   �   �          %          m_valid => dv      ( j   ),�   �   �          $          m_dataZ => wirez   ( j+1 )�   �   �          %          m_dataY => wirey   ( j+1 ),�   �   �          %          m_dataX => wirex   ( j+1 ),5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n�     �   �   �   �      +                 m_dataZ => wirez   ( j+1 )5�_�  �  �          �   �       ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n�     �   �   �   �                     rst     => rst,5�_�  �  �          �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n�     �   �   �                      );�   �   �                         rst     => rst�   �   �                         clk     => clk,�   �   �                      s_atan  =>�   �   �          '            s_inv   => inv     ( j   ),�   �   �          '            s_ready => en      ( j   ),�   �   �                   s_valid =>�   �   �          $         s_dataT => wireLUT ( j   ),�   �   �          $         s_dataZ => wirez   ( j   ),�   �   �          $         s_dataY => wirey   ( j   ),�   �   �          $         s_dataX => wirex   ( j   ),�   �   �                m_ready =>�   �   �          !      m_inv   => inv     ( j+1 ),�   �   �          !      m_valid => dv      ( j   ),5�_�  �     �      �   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   �   �   �                       m_ready =>5�_�  �                @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');5�_�                  @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   ?   A   �      H   signal en, dv, inv, rdy            : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   ?   A   �      G   signal en, dv, inv, rdy           : handShakeVector:= (others=>'0');5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   �   �   �                       m_ready => 5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^n�     �   �   �   �                          s_valid =>5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o     �   �   �   �    �   �   �   �    5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o     �   ?   A   �      F   signal en, dv, inv, rdy          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o     �   ?   A   �      H   signal en, dv, inv, s_rdy          : handShakeVector:= (others=>'0');5�_�    	             @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o     �   ?   A   �      P   signal en, dv, inv, s_rdy,m_valid          : handShakeVector:= (others=>'0');5�_�    
          	   �   	    ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o(     �   �   �   �               en(j+1)<=dv(j);5�_�  	            
   �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o+     �   �   �   �               s_rdyen(j+1)<=dv(j);5�_�  
               �       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o+     �   �   �   �               s_rdyn(j+1)<=dv(j);5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      Q   signal en, dv, inv, s_rdy, m_valid          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      R   signal en, dv, inv, s_rdy, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      S   signal en, dv, inv, sw_rdy, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      V   signal en, dv, inv, sw_readdy, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      U   signal en, dv, inv, sw_ready, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @       ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      T   signal en, dv, inv, s_ready, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @   "    ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      U   signal en, dv, inv, s_readyW, mw_valid          : handShakeVector:= (others=>'0');5�_�                 @   (    ����                                                                                                                                                                                                                                                                                                                            �           �           V        ^o�     �   ?   A   �      T   signal en, dv, inv, s_readyW, m_valid          : handShakeVector:= (others=>'0');5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �          �   !       v   !    ^o�     �   �   �   �      "                    s_valid => rdy�   �   �   �    5�_�                 �   -    ����                                                                                                                                                                                                                                                                                                                            �          �   -       v   !    ^o�     �   �   �   �    5�_�                 �        ����                                                                                                                                                                                                                                                                                                                            �          �   -       v   !    ^o�     �   �   �           5�_�                 �   "    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^o�     �   �   �   �      2                       s_ready => en      ( j   ),5�_�                 �   "    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p     �   �   �   �      #                       s_ready => ,5�_�                 �   $    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p	     �   �   �   �      %                       s_ready => m_,5�_�                 �   )    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p     �   �   �   �      +                       s_ready => m_valid(,5�_�                 �   +    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �      ,                       s_ready => m_validW(,5�_�                 �   	    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �               s_rdy(j+1)<=dv(j);5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �               m_validW(j+1)<=dv(j);5�_�                 �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �               m_validW(j1)<=dv(j);5�_�                  �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �               m_validW(j)<=dv(j);5�_�    !              �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �               m_validW(j+1)<=dv(j);5�_�     "          !   �   "    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �      .                       s_ready => m_validW(j),5�_�  !  #          "   �   	    ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �      $         m_validW(j+1)<=s_readyW(j);5�_�  "  $          #   �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �      $         s_readyW(j+1)<=s_readyW(j);5�_�  #  %          $   �       ����                                                                                                                                                                                                                                                                                                                            �   "       �   0       v   0    ^p�     �   �   �   �      $         s_readyW(j+1)<=m_readyW(j);5�_�  $  &          %   �       ����                                                                                                                                                                                                                                                                                                                            �          �          v       ^q     �   �   �   �      $         s_readyW(j+1)<=m_readyW(j);5�_�  %  (          &   �        ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^q     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_validW(j);�   �   �   �                en(j+1)       <= dv(j);�   �   �   �                             );�   �   �   �      (                          rst     => rst�   �   �   �      )                          clk     => clk,�   �   �   �      !                       s_atan  =>�   �   �   �      2                       s_inv   => inv     ( j   ),�   �   �   �      .                       s_ready => s_readyW(j),�   �   �   �      .                    s_valid => en      ( j   )�   �   �   �      /                    s_dataT => wireLUT ( j   ),�   �   �   �      /                    s_dataZ => wirez   ( j   ),�   �   �   �      /                    s_dataY => wirey   ( j   ),�   �   �   �      /                    s_dataX => wirex   ( j   ),�   �   �   �      !                 m_ready => rdy (�   �   �   �      ,                 m_inv   => inv     ( j+1 ),�   �   �   �      ,                 m_valid => dv      ( j   ),�   �   �   �      ,                 m_dataZ => wirez   ( j+1 ),�   �   �   �      ,                 m_dataY => wirey   ( j+1 ),�   �   �   �      ,                 m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      !                  en ( 0 )<= '0';�   w   y   �      $               when waitingCordic =>�   v   x   �                        end if;�   u   w   �      2                     bitCounter := bitCounter + 1;�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      @                          state                <= waitingCordic;�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   n   p   �      !                          end if;�   m   o   �      :                                wirez(0) <= (others=>'0');�   l   n   �                                else �   k   m   �      $                             end if;�   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   i   k   �      "                             else �   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   g   i   �      8                             if s_axis_tdata(7)='1' then�   f   h   �      ,                          if inv(0)='1' then�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   d   f   �      4                          wirey(0) <= (others=>'0');�   c   e   �      !                        when 1 =>�   b   d   �      !                          end if;�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   [   ]   �      4                          wirex(0) <= (others=>'0');�   Z   \   �      !                        when 0 =>�   Y   [   �      '                     case bitCounter is�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case state is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      U   signal en, dv, inv, s_readyW, m_validW          : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                   en(j+1)<=dv(j);�   �   �          $         s_readyW(j+1)<=m_validW(j);5�_�  &  )  '      (   T        ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^q7     �   S   U   �    �   T   U   �    5�_�  (  *          )   U       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^qi     �   T   V   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada5�_�  )  +          *   U       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^qn     �   T   V   �      Y            s_readyW(0)        <= '0';                           --y ya no tengo mas nada5�_�  *  ,          +   U   !    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^qq     �   T   V   �      T            s_readyW(0)   <= '0';                           --y ya no tengo mas nada5�_�  +  -          ,   �       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^r
     �   �   �   �      &         s_readyW(j+1) <= m_validW(j);5�_�  ,  .          -   @   #    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^r     �   ?   A   �      U   signal en, dv, inv, s_readyW, m_validW          : handShakeVector:= (others=>'0');5�_�  -  /          .   @   !    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   ?   A   �      U   signal en, dv, inv, s_readyW, m_readyW          : handShakeVector:= (others=>'0');5�_�  .  0          /   �       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      !                 m_ready => rdy (5�_�  /  1          0   �   $    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      )                 m_ready => m_readyWrdy (5�_�  0  2          1   �   &    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      +                 m_ready => m_readyW(jrdy (5�_�  1  3          2   �   &    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      &                 m_ready => m_readyW(j5�_�  2  4          3   �   '    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      '                 m_ready => m_readyW(j)5�_�  3  5          4   �   '    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^s�     �   �   �   �      (                 m_ready => m_readyW(j)m5�_�  4  6          5   @   
    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t     �   ?   A   �      U   signal en, dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  5  7          6   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t     �   ?   A   �      \   signal s_validen, dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  6  8          7   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t     �   ?   A   �      ]   signal s_validWen, dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  7  9          8   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t     �   ?   A   �      \   signal s_validWe, dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  8  :          9   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t     �   ?   A   �      [   signal s_validW, dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  9  ;          :   @   )    ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t'     �   ?   A   �      ]   signal s_validW, s_dv, inv, s_readyW, s_readyW          : handShakeVector:= (others=>'0');5�_�  :  <          ;   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t*     �   ?   A   �      ]   signal s_validW, s_dv, inv, s_readyW, m_readyW          : handShakeVector:= (others=>'0');5�_�  ;  =          <   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t+     �   ?   A   �      ]   signal s_validW, m_dv, inv, s_readyW, m_readyW          : handShakeVector:= (others=>'0');5�_�  <  >          =   @       ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^t,     �   ?   A   �      \   signal s_validW, m_v, inv, s_readyW, m_readyW          : handShakeVector:= (others=>'0');5�_�  =  ?          >   @       ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t0     �   ?   A   �      a   signal s_validW, m_validW, inv, s_readyW, m_readyW          : handShakeVector:= (others=>'0');5�_�  >  @          ?   @   /    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t2     �   ?   A   �      \   signal s_validW, m_validW, s_readyW, m_readyW          : handShakeVector:= (others=>'0');�   @   A   �    5�_�  ?  A          @   @   0    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t5     �   ?   A   �      a   signal s_validW, m_validW, s_readyW, m_readyWinv,           : handShakeVector:= (others=>'0');5�_�  @  B          A   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t7     �   ?   A   �      b   signal s_validW, m_validW, s_readyW, m_readyW,inv,           : handShakeVector:= (others=>'0');5�_�  A  C          B   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t7     �   ?   A   �      a   signal s_validW, m_validW, s_readyW, m_readyW,inv           : handShakeVector:= (others=>'0');5�_�  B  D          C   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t7     �   ?   A   �      `   signal s_validW, m_validW, s_readyW, m_readyW,inv          : handShakeVector:= (others=>'0');5�_�  C  E          D   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t7     �   ?   A   �      _   signal s_validW, m_validW, s_readyW, m_readyW,inv         : handShakeVector:= (others=>'0');5�_�  D  F          E   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t7     �   ?   A   �      ^   signal s_validW, m_validW, s_readyW, m_readyW,inv        : handShakeVector:= (others=>'0');5�_�  E  G          F   @   4    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t8     �   ?   A   �      ]   signal s_validW, m_validW, s_readyW, m_readyW,inv       : handShakeVector:= (others=>'0');5�_�  F  H          G   @   6    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^t9     �   ?   A   �      \   signal s_validW, m_validW, s_readyW, m_readyW,inv      : handShakeVector:= (others=>'0');5�_�  G  I          H   S       ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^tB     �   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada5�_�  H  J          I   q       ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^tV     �   p   r   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada5�_�  I  K          J   q   !    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^tj     �   p   r   �      n                          s_valid(0)                <= '1';                           --y ya no tengo mas nada5�_�  J  L          K   q   "    ����                                                                                                                                                                                                                                                                                                                            @          @   "       v   "    ^tk     �   p   r   �      p                          s_validWE(0)                <= '1';                           --y ya no tengo mas nada5�_�  K  M          L   q        ����                                                                                                                                                                                                                                                                                                                            q   ,       t   ,       V   ,    ^to     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �                en(j+1)       <= dv(j);�   �   �   �                             );�   �   �   �      (                          rst     => rst�   �   �   �      )                          clk     => clk,�   �   �   �      !                       s_atan  =>�   �   �   �      2                       s_inv   => inv     ( j   ),�   �   �   �      .                       s_ready => s_readyW(j),�   �   �   �      .                    s_valid => en      ( j   )�   �   �   �      /                    s_dataT => wireLUT ( j   ),�   �   �   �      /                    s_dataZ => wirez   ( j   ),�   �   �   �      /                    s_dataY => wirey   ( j   ),�   �   �   �      /                    s_dataX => wirex   ( j   ),�   �   �   �      (                 m_ready => m_readyW(j),�   �   �   �      ,                 m_inv   => inv     ( j+1 ),�   �   �   �      ,                 m_valid => dv      ( j   ),�   �   �   �      ,                 m_dataZ => wirez   ( j+1 ),�   �   �   �      ,                 m_dataY => wirey   ( j+1 ),�   �   �   �      ,                 m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   p   r          o                          s_validW(0)                <= '1';                           --y ya no tengo mas nada�   s   u          @                          state                <= waitingCordic;�   r   t          i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   q   s          r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo5�_�  L  N          M   �       ����                                                                                                                                                                                                                                                                                                                            q   ,       t   ,       V   ,    ^t     �   �   �   �      .                    s_valid => en      ( j   )5�_�  M  O          N   �   '    ����                                                                                                                                                                                                                                                                                                                            q   ,       t   ,       V   ,    ^t�     �   �   �   �      4                    s_valid => s_validW      ( j   )5�_�  N  P          O           ����                                                                                                                                                                                                                                                                                                                            q   ,       t   ,       V   ,    ^t�     �          �      library IEEE;5�_�  O  Q          P   {       ����                                                                                                                                                                                                                                                                                                                            q   ,       t   ,       V   ,    ^t�     �   z   |   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo5�_�  P  R          Q   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^t�     �   �   �   �      ,                 m_valid => dv      ( j   ),5�_�  Q  S          R   �   $    ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^t�     �   �   �   �      2                 m_valid => m_validW      ( j   ),5�_�  R  T          S   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^t�     �   �   �   �                en(j+1)       <= dv(j);5�_�  S  U          T   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^t�     �   �   �   �               en(j+1)       <= (j);5�_�  T  V          U   �   	    ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^t�     �   �   �   �      &         en(j+1)       <= m_validW(j);5�_�  U  W          V   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t�     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �                             );�   �   �   �      (                          rst     => rst�   �   �   �      )                          clk     => clk,�   �   �   �      !                       s_atan  =>�   �   �   �      2                       s_inv   => inv     ( j   ),�   �   �   �      .                       s_ready => s_readyW(j),�   �   �   �      .                    s_valid => s_validW( j   )�   �   �   �      /                    s_dataT => wireLUT ( j   ),�   �   �   �      /                    s_dataZ => wirez   ( j   ),�   �   �   �      /                    s_dataY => wirey   ( j   ),�   �   �   �      /                    s_dataX => wirex   ( j   ),�   �   �   �      (                 m_ready => m_readyW(j),�   �   �   �      ,                 m_inv   => inv     ( j+1 ),�   �   �   �      ,                 m_valid => m_validW( j   ),�   �   �   �      ,                 m_dataZ => wirez   ( j+1 ),�   �   �   �      ,                 m_dataY => wirey   ( j+1 ),�   �   �   �      ,                 m_dataX => wirex   ( j+1 ),�   �   �   �            port map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          ,         s_validW(j+1)       <= m_validW(j);�   �   �          &         s_readyW(j+1) <= m_readyW(j);5�_�  V  X          W   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t�     �   �   �          !                       s_atan  =>5�_�  W  Y          X   �        ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �                                 );�   �   �          (                          rst     => rst�   �   �          )                          clk     => clk,�   �   �          2                       s_inv   => inv     ( j   ),�   �   �          .                       s_ready => s_readyW(j),�   �   �          .                    s_valid => s_validW( j   )�   �   �          /                    s_dataT => wireLUT ( j   ),�   �   �          /                    s_dataZ => wirez   ( j   ),�   �   �          /                    s_dataY => wirey   ( j   ),�   �   �          /                    s_dataX => wirex   ( j   ),5�_�  X  Z          Y   �   +    ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �   �      +                 s_valid => s_validW( j   )5�_�  Y  [          Z   �   +    ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �   �      ,                 s_valid => s_validW( j   )m5�_�  Z  \          [   �        ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �             );�   �   �                rst     => rst�   �   �                clk     => clk,�   �   �          !      s_inv   => inv     ( j   ),�   �   �                s_ready => s_readyW(j),5�_�  [  ]          \   �        ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �                    );�   �   �   �                       rst     => rst�   �   �   �                        clk     => clk,�   �   �   �      .                 s_inv   => inv       ( j   ),�   �   �   �      (                 s_ready => s_readyW(j),�   �   �   �      *                 s_valid => s_validW( j ),�   �   �   �      .                 s_dataT => wireLUT   ( j   ),�   �   �   �      .                 s_dataZ => wirez     ( j   ),�   �   �   �      .                 s_dataY => wirey     ( j   ),�   �   �   �      .                 s_dataX => wirex     ( j   ),�   �   �   �      (                 m_ready => m_readyW(j),�   �   �   �      .                 m_inv   => inv       ( j+1 ),�   �   �   �      *                 m_valid => m_validW( j ),�   �   �   �      .                 m_dataZ => wirez     ( j+1 ),�   �   �   �      .                 m_dataY => wirey     ( j+1 ),�   �   �   �      .                 m_dataX => wirex     ( j+1 ),�   �   �   �            port               map(�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                           rst     => rst�   �   �                            clk     => clk,�   �   �          ,                 s_inv   => inv     ( j   ),�   �   �          (                 s_ready => s_readyW(j),�   �   �          ,                 s_valid => s_validW( j   ),�   �   �          ,                 s_dataT => wireLUT ( j   ),�   �   �          ,                 s_dataZ => wirez   ( j   ),�   �   �          ,                 s_dataY => wirey   ( j   ),�   �   �          ,                 s_dataX => wirex   ( j   ),�   �   �          (                 m_ready => m_readyW(j),�   �   �          ,                 m_inv   => inv     ( j+1 ),�   �   �          ,                 m_valid => m_validW( j   ),�   �   �          ,                 m_dataZ => wirez   ( j+1 ),�   �   �          ,                 m_dataY => wirey   ( j+1 ),�   �   �          ,                 m_dataX => wirex   ( j+1 ),�   �   �                port map(5�_�  \  ^          ]   �       ����                                                                                                                                                                                                                            �                                                                                              �           �          V       ^t�     �   �   �   �            port               map(5�_�  ]  _          ^   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t�     �   �   �   �      .                 m_dataX => wirex     ( j+1 ),   .                 m_dataY => wirey     ( j+1 ),   .                 m_dataZ => wirez     ( j+1 ),   *                 m_valid => m_validW( j ),   .                 m_inv   => inv       ( j+1 ),   (                 m_ready => m_readyW(j),       .                 s_dataX => wirex     ( j   ),   .                 s_dataY => wirey     ( j   ),   .                 s_dataZ => wirez     ( j   ),   .                 s_dataT => wireLUT   ( j   ),   *                 s_valid => s_validW( j ),   (                 s_ready => s_readyW(j),   .                 s_inv   => inv       ( j   ),                         clk     => clk,                    rst     => rst5�_�  ^  `          _   �        ����                                                                                                                                                                                                                            �                                                                                              �          �           v        ^t�     �   �   �                  rst     => rst�   �   �                  clk     => clk,�   �   �          %        s_inv   => inv       ( j   ),�   �   �                  s_ready => s_readyW(j),�   �   �          !        s_valid => s_validW( j ),�   �   �          %        s_dataT => wireLUT   ( j   ),�   �   �          %        s_dataZ => wirez     ( j   ),�   �   �          %        s_dataY => wirey     ( j   ),�   �   �          %        s_dataX => wirex     ( j   ),�   �   �                  m_ready => m_readyW(j),�   �   �          %        m_inv   => inv       ( j+1 ),�   �   �          !        m_valid => m_validW( j ),�   �   �          %        m_dataZ => wirez     ( j+1 ),�   �   �          %        m_dataY => wirey     ( j+1 ),�   �   �          %        m_dataX => wirex     ( j+1 ),5�_�  _  a          `   �        ����                                                                                                                                                                                                                            �                                                                                              �          �           v        ^t�     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �      -                                           );�   �   �   �                       rst     => rst�   �   �   �                        clk     => clk,�   �   �   �      -                 s_inv   => inv      ( j   ),�   �   �   �      -                 s_ready => s_readyW ( j   ),�   �   �   �      -                 s_valid => s_validW ( j   ),�   �   �   �      -                 s_dataT => wireLUT  ( j   ),�   �   �   �      -                 s_dataZ => wirez    ( j   ),�   �   �   �      -                 s_dataY => wirey    ( j   ),�   �   �   �      -                 s_dataX => wirex    ( j   ),�   �   �   �      -                 m_ready => m_readyW ( j   ),�   �   �   �      -                 m_inv   => inv      ( j+1 ),�   �   �   �      -                 m_valid => m_validW ( j   ),�   �   �   �      -                 m_dataZ => wirez    ( j+1 ),�   �   �   �      -                 m_dataY => wirey    ( j+1 ),�   �   �   �      -                 m_dataX => wirex    ( j+1 ),�   �   �   �      &      port map                       (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                        );�   �   �          +                 s_valid => s_validW ( j ),�   �   �          -                 s_dataT => wireLUT  ( j   ),�   �   �          -                 m_inv   => inv      ( j+1 ),�   �   �          -                 s_dataY => wirey    ( j   ),�   �   �          -                 m_dataZ => wirez    ( j+1 ),�   �   �          -                 m_dataY => wirey    ( j+1 ),�   �   �          *                 s_ready => s_readyW ( j),�   �   �          -                 m_dataX => wirex    ( j+1 ),�   �   �          *                 m_ready => m_readyW ( j),�   �   �          +                 m_valid => m_validW ( j ),�   �   �          -                 s_dataZ => wirez    ( j   ),�   �   �          -                 s_inv   => inv      ( j   ),�   �   �          -                 s_dataX => wirex    ( j   ),�   �   �          *                 s_valid => s_validW( j ),�   �   �          .                 s_dataT => wireLUT   ( j   ),�   �   �          .                 m_inv   => inv       ( j+1 ),�   �   �          .                 s_dataY => wirey     ( j   ),�   �   �          .                 m_dataZ => wirez     ( j+1 ),�   �   �          .                 m_dataY => wirey     ( j+1 ),�   �   �          (                 s_ready => s_readyW(j),�   �   �                port map(�   �   �          .                 m_dataX => wirex     ( j+1 ),�   �   �          (                 m_ready => m_readyW(j),�   �   �          *                 m_valid => m_validW( j ),�   �   �          .                 s_dataZ => wirez     ( j   ),�   �   �          .                 s_inv   => inv       ( j   ),�   �   �          .                 s_dataX => wirex     ( j   ),5�_�  `  b          a   �        ����                                                                                                                                                                                                                            �                                                                                              �          �           v        ^t�     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �      -                                           );�   �   �   �                        rst     =>  rst�   �   �   �      !                 clk     =>  clk,�   �   �   �      .                 s_inv   =>  inv      ( j   ),�   �   �   �      .                 s_ready =>  s_readyW ( j   ),�   �   �   �      .                 s_valid =>  s_validW ( j   ),�   �   �   �      .                 s_dataT =>  wireLUT  ( j   ),�   �   �   �      .                 s_dataZ =>  wirez    ( j   ),�   �   �   �      .                 s_dataY =>  wirey    ( j   ),�   �   �   �      .                 s_dataX =>  wirex    ( j   ),�   �   �   �      .                 m_ready =>  m_readyW ( j   ),�   �   �   �      .                 m_inv   =>  inv      ( j+1 ),�   �   �   �      .                 m_valid =>  m_validW ( j   ),�   �   �   �      .                 m_dataZ =>  wirez    ( j+1 ),�   �   �   �      .                 m_dataY =>  wirey    ( j+1 ),�   �   �   �      .                 m_dataX =>  wirex    ( j+1 ),�   �   �   �            port               map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                           rst     => rst�   �   �                            clk     => clk,�   �   �          -                 s_inv   => inv      ( j   ),�   �   �          -                 s_ready => s_readyW ( j   ),�   �   �          -                 s_valid => s_validW ( j   ),�   �   �          -                 s_dataT => wireLUT  ( j   ),�   �   �          -                 s_dataZ => wirez    ( j   ),�   �   �          -                 s_dataY => wirey    ( j   ),�   �   �          -                 s_dataX => wirex    ( j   ),�   �   �          -                 m_ready => m_readyW ( j   ),�   �   �          -                 m_inv   => inv      ( j+1 ),�   �   �          -                 m_valid => m_validW ( j   ),�   �   �          -                 m_dataZ => wirez    ( j+1 ),�   �   �          -                 m_dataY => wirey    ( j+1 ),�   �   �          -                 m_dataX => wirex    ( j+1 ),�   �   �          &      port map                       (5�_�  a  c          b   �        ����                                                                                                                                                                                                                            �                                                                                              �          �           v        ^t�     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �      -                                           );�   �   �   �                       rst     => rst�   �   �   �                        clk     => clk,�   �   �   �      -                 s_inv   => inv      ( j   ),�   �   �   �      -                 s_ready => s_readyW ( j   ),�   �   �   �      -                 s_valid => s_validW ( j   ),�   �   �   �      -                 s_dataT => wireLUT  ( j   ),�   �   �   �      -                 s_dataZ => wirez    ( j   ),�   �   �   �      -                 s_dataY => wirey    ( j   ),�   �   �   �      -                 s_dataX => wirex    ( j   ),�   �   �   �      -                 m_ready => m_readyW ( j   ),�   �   �   �      -                 m_inv   => inv      ( j+1 ),�   �   �   �      -                 m_valid => m_validW ( j   ),�   �   �   �      -                 m_dataZ => wirez    ( j+1 ),�   �   �   �      -                 m_dataY => wirey    ( j+1 ),�   �   �   �      -                 m_dataX => wirex    ( j+1 ),�   �   �   �            port               map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�      �   �                        end if;�   ~   �   �      (                     bitCounter    := 0;�   }      �      4                     state         <= waitingMready;�   |   ~   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   {   }   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   z   |   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   y   {   �      !                  en ( 0 )<= '0';�   x   z   �      $               when waitingCordic =>�   w   y   �                        end if;�   v   x   �      2                     bitCounter := bitCounter + 1;�   u   w   �                           end case;�   t   v   �      &                        when others =>�   s   u   �      9                          state         <= waitingCordic;�   r   t   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   q   s   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   p   r   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   o   q   �      !                          end if;�   n   p   �      :                                wirez(0) <= (others=>'0');�   m   o   �                                else �   l   n   �      $                             end if;�   k   m   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   j   l   �      "                             else �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   h   j   �      8                             if s_axis_tdata(7)='1' then�   g   i   �      ,                          if inv(0)='1' then�   f   h   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   e   g   �      4                          wirey(0) <= (others=>'0');�   d   f   �      !                        when 1 =>�   c   e   �      !                          end if;�   b   d   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   a   c   �      -                             inv(0)   <= '0';�   `   b   �                                else�   _   a   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '1';�   ]   _   �      5                          if s_axis_tdata(7)='1' then�   \   ^   �      4                          wirex(0) <= (others=>'0');�   [   ]   �      !                        when 0 =>�   Z   \   �      '                     case bitCounter is�   Y   [   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   X   Z   �      $               when waitingSvalid =>�   W   Y   �                  case state is�   V   X   �               else�   U   W   �                  bitCounter    := 0;�   T   V   �      !            s_readyW(0)   <= '0';�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   R   T   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   Q   S   �      -            angle         <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   N   P   �      !            m_axis_tvalid <= '0';�   M   O   �      !            s_axis_tready <= '1';�   L   N   �      +            state         <= waitingSvalid;�   K   M   �               if rst = '0' then�   J   L   �            if rising_edge(clk) then�   I   K   �         begin�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   G   I   �      *      variable sign :signed (15 downto 0);�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �      %   cordic_proc:process (clk) is --{{{�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �         �   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   8   :   �      '   signal clockWise : std_logic := '0';�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �         end component; --}}}�   0   2   �                );�   /   1   �      )          rst           : in  STD_LOGIC);�   .   0   �      (          clk           : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �                            rst     =>  rst�   �   �          !                 clk     =>  clk,�   �   �          .                 s_inv   =>  inv      ( j   ),�   �   �          .                 s_ready =>  s_readyW ( j   ),�   �   �          .                 s_valid =>  s_validW ( j   ),�   �   �          .                 s_dataT =>  wireLUT  ( j   ),�   �   �          .                 s_dataZ =>  wirez    ( j   ),�   �   �          .                 s_dataY =>  wirey    ( j   ),�   �   �          .                 s_dataX =>  wirex    ( j   ),�   �   �          .                 m_ready =>  m_readyW ( j   ),�   �   �          .                 m_inv   =>  inv      ( j+1 ),�   �   �          .                 m_valid =>  m_validW ( j   ),�   �   �          .                 m_dataZ =>  wirez    ( j+1 ),�   �   �          .                 m_dataY =>  wirey    ( j+1 ),�   �   �          .                 m_dataX =>  wirex    ( j+1 ),5�_�  b  d          c   �       ����                                                                                                                                                                                                                            �                                                                                              �          �           v        ^t�     �   �   �   �            port               map (5�_�  c  e          d   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t�     �   �   �   �      -                 m_dataX => wirex    ( j+1 ),   -                 m_dataY => wirey    ( j+1 ),   -                 m_dataZ => wirez    ( j+1 ),   -                 m_valid => m_validW ( j   ),   -                 m_inv   => inv      ( j+1 ),   -                 m_ready => m_readyW ( j   ),       -                 s_dataX => wirex    ( j   ),   -                 s_dataY => wirey    ( j   ),   -                 s_dataZ => wirez    ( j   ),   -                 s_dataT => wireLUT  ( j   ),   -                 s_valid => s_validW ( j   ),   -                 s_ready => s_readyW ( j   ),   -                 s_inv   => inv      ( j   ),                         clk     => clk,                    rst     => rst5�_�  d  f          e   �   	    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t�    �   �   �   �      -                                           );5�_�  e  g          f   ;        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u   �   :   <   �         5�_�  f  h          g           ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u   �          �      IEEE;5�_�  g  i          h   1   
    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u   �   0   1                    );5�_�  h  j          i           ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u)   �          �      	use IEEE;5�_�  i  k          j   y       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u1     �   x   z   �      !                  en ( 0 )<= '0';5�_�  j  l          k   y       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^uP     �   x   z   �      '                  s_valide ( 0 )<= '0';5�_�  k  m          l   y       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^uP   �   x   z   �      (                  s_validWe ( 0 )<= '0';5�_�  l  n          m   -        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u�   �   ,   -          "          s_atan  : in  STD_LOGIC;5�_�  m  o          n   x        ����                                                                                                                                                                                                                            �                                                                                              x   &       x   &       V   *    ^��     �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => s_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j   ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => m_validW ( j   ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�      �   �      $               when waitingMready =>�   }      �                        end if;�   |   ~   �      (                     bitCounter    := 0;�   {   }   �      4                     state         <= waitingMready;�   z   |   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   y   {   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   x   z   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   w   y   �      (                  s_validW ( 0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            s_readyW(0)   <= '0';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   w   y          '                  s_validW ( 0 )<= '0';5�_�  n  p          o   K        ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��   �   �   �   �         end generate;�   �   �   �      &         s_readyW(j+1) <= m_readyW(j);�   �   �   �      &         s_validW(j+1) <= m_validW(j);�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => s_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j   ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => m_validW ( j   ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�      �   �      $               when waitingMready =>�   }      �                        end if;�   |   ~   �      (                     bitCounter    := 0;�   {   }   �      4                     state         <= waitingMready;�   z   |   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   y   {   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   x   z   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo�   w   y   �      (                  s_validW ( 0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            s_readyW(0)   <= '0';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            s_validW(0)   <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   J   L          +            state         <= waitingSvalid;�   N   P          !            clockWise     <= '0';�   S   U                      bitCounter    := 0;�   R   T          !            s_readyW(0)   <= '0';�   L   N          !            m_axis_tvalid <= '0';�   P   R          Z            s_validW(0)         <= '0';                           --y ya no tengo mas nada�   O   Q          -            angle         <= (others => '0');�   K   M          !            s_axis_tready <= '1';�   Q   S          T            inv(0)        <= '0';                           --y ya no tengo mas nada�   M   O          -            m_axis_tdata  <= (others => '0');5�_�  o  q          p   S       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�N   �   R   T   �      !            s_readyW(0)   <= '0';5�_�  p  r          q   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      '           s_ready => s_readyW ( j   ),5�_�  q  s          r   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      '           s_ready => m_readyW ( j   ),5�_�  r  t          s   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�/     �   �   �   �      '           m_ready => m_readyW ( j   ),5�_�  s  u          t   �   "    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�1     �   �   �   �      '           m_ready => s_readyW ( j   ),5�_�  t  v          u   �   $    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�2     �   �   �   �      )           m_ready => s_readyW ( j+1   ),5�_�  u  w          v   �   $    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�3     �   �   �   �      (           m_ready => s_readyW ( j+1  ),5�_�  v  x          w   �        ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      &         s_readyW(j+1) <= m_readyW(j);5�_�  w  y          x   �        ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      (00         s_readyW(j+1) <= m_readyW(j);5�_�  x  z          y   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      '           m_ready => s_readyW ( j+1 ),5�_�  y  {          z   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   �   �   �      '           m_ready => n_readyW ( j+1 ),5�_�  z  |          {   �       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��  	 �   �   �   �      '           m_ready => n_readyW ( j+1 ),5�_�  {  }          |   S       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�     �   R   T   �      !            s_readyW(0)   <= '1';5�_�  |  ~          }   S       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�  
 �   R   T   �      !            m_readyW(0)   <= '1';5�_�  }            ~   o   /    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�     �   n   p   �      G                          s_validW(0)   <= '1';--y ya no tengo mas nada5�_�  ~  �             y       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^�L     �   x   z   �      p                  if m_validW(0) = '1' then                           --espero e que este listo para enviar algo5�_�    �          �   y       ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   x   z   �      p                  if m_readyW(0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   y   "    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   x   z   �      u                  if m_readyW(ITER-1) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �  �      �   y   "    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��   �   x   z   �      t                  if m_readyW(ITER1) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �  �      �   y       ����                                                                                                                                                                                                                            �                                                                                              y          ~                 ^�w     �   x   z   �    �   y   z   �    5�_�  �  �          �   z       ����                                                                                                                                                                                                                            �                                                                                              z                           ^�z   �   z   �   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);   ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada   4                     state         <= waitingMready;   (                     bitCounter    := 0;                     end if;�   y   {   �      s                  if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�z   �   w   y   �      (                  s_validW ( 0 ) <= '0';5�_�  �  �          �   �   "    ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   �   �   �      '           m_valid => m_validW ( j   ),5�_�  �  �          �   �   $    ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   �   �   �      *           m_valid => m_validW ( j+1l   ),5�_�  �  �          �   �   $    ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   �   �   �      )           m_valid => m_validW ( j+1   ),5�_�  �  �          �   �   $    ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   �   �   �      (           m_valid => m_validW ( j+1  ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   �   �   �      '           m_valid => m_validW ( j+1 ),5�_�  �  �          �   �        ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�'     �   �   �   �      &         s_validW(j+1) <= m_validW(j);5�_�  �  �          �   �        ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�)     �   �   �   �      (00         s_validW(j+1) <= m_validW(j);5�_�  �  �          �   �        ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�,     �   �   �   �      (00R        s_validW(j+1) <= m_validW(j);5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�.     �   �   �   �      (--R        s_validW(j+1) <= m_validW(j);5�_�  �  �          �   >       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >          v       ^�4   �   =   ?   �      X   signal s_validW, m_validW, s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >          v       ^��     �   w   y   �      *                  --s_validW ( 0 ) <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >          v       ^��   �   w   y   �      )                  -s_validW ( 0 ) <= '0';5�_�  �  �          �   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          '--        s_validW(j+1) <= m_validW(j);   (--         s_readyW(j+1) <= m_readyW(j);5�_�  �  �          �   >   
    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   =   ?   �      O   signal s_validW,  s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   >   
    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   =   ?   �      N   signal _validW,  s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   >       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   =   ?   �      M   signal validW,  s_readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   >       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   =   ?   �      L   signal validW,  _readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   >       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��   �   =   ?   �      K   signal validW,  readyW, m_readyW,inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   Q       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   P   R   �      T            s_validW(0)   <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   Q       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   P   R   �      S            _validW(0)   <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   Q       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��   �   P   R   �      R            validW(0)   <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   S       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   R   T   �      !            m_readyW(0)   <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   R   T   �                   _readyW(0)   <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��   �   R   T   �                  readyW(0)   <= '1';5�_�  �  �          �   o       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   n   p   �      /                          s_validW(0)   <= '1';5�_�  �  �          �   o       ����                                                                                                                                                                >   
                                                       �                                                                                              >          >   "       v   "    ^��     �   n   p   �      .                          _validW(0)   <= '1';5�_�  �  �          �   o        ����                                                                                                                                                                >   
                                                       �                                                                                              o          r          V       ^��     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y   �      (                  s_validW ( 0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   n   p          -                          validW(0)   <= '1';�   q   s          9                          state         <= waitingCordic;�   p   r          b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q          k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              o          r          V       ^�     �   w   y   �      (                  s_validW ( 0 ) <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              o          r          V       ^�     �   w   y   �      '                  _validW ( 0 ) <= '0';5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�   �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y   �      *                  validW ( 0 )     <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   w   y          &                  validW ( 0 ) <= '0';�   x   z          ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y   �      1                  validW           (  0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   x   z          ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y          *                  validW ( 0 )     <= '0';5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�
     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      d                     m_axis_tvalid        <= '1';                           --y ya no tengo mas nada�   w   y   �      1                  validW           (  0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   w   y          1                  validW           (  0 ) <= '0';�   x   z          ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   y        ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   x   z          d                     m_axis_tvalid        <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x   "       y   "       V   "    ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      Z                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y   �      .                  validW        (  0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   x   z          a                  m_axis_tvalid        <= '1';                           --y ya no tengo mas nada�   w   y          1                  validW           (  0 ) <= '0';5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      a                  m_axis_tvalid        <= '1';                           --y ya no tengo mas nada�   w   y   �      .                  validW        (  0 ) <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   w   y          .                  validW        (  0 ) <= '0';�   x   z          Z                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   w   y   �      .                  validW        (  0 ) <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   w   y   �      -                  validW       (  0 ) <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   w   y   �      &                  validW(  0 ) <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x           y           V        ^�     �   w   y   �      $                  validW(0 ) <= '0';5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�   �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => m_readyW ( j   ),�   �   �   �      '           s_valid => s_validW ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => m_readyW ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => s_validW ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        --end if;�   }      �      *                  --   bitCounter    := 0;�   |   ~   �      6                  --   state         <= waitingMready;�   {   }   �      _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      Z                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   w   y   �      '                  validW(0)     <= '0';�   v   x   �      $               when waitingCordic =>�   u   w   �                        end if;�   t   v   �      2                     bitCounter := bitCounter + 1;�   s   u   �                           end case;�   r   t   �      &                        when others =>�   q   s   �      9                          state         <= waitingCordic;�   p   r   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   o   q   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      :                                wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      ,                          if inv(0)='1' then�   d   f   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   c   e   �      4                          wirey(0) <= (others=>'0');�   b   d   �      !                        when 1 =>�   a   c   �      !                          end if;�   `   b   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   _   a   �      -                             inv(0)   <= '0';�   ^   `   �                                else�   ]   _   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   \   ^   �      -                             inv(0)   <= '1';�   [   ]   �      5                          if s_axis_tdata(7)='1' then�   Z   \   �      4                          wirex(0) <= (others=>'0');�   Y   [   �      !                        when 0 =>�   X   Z   �      '                     case bitCounter is�   W   Y   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   V   X   �      $               when waitingSvalid =>�   U   W   �                  case state is�   T   V   �               else�   S   U   �                  bitCounter    := 0;�   R   T   �      !            readyW(0)     <= '1';�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   w   y          #                  validW(0) <= '0';�   x   z          a                  m_axis_tvalid        <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�$     �   �   �   �      '           m_valid => s_validW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�$     �   �   �   �      &           m_valid => _validW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�&     �   �   �   �      %           m_valid => validW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�)     �   �   �   �      '           s_valid => s_validW ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�)     �   �   �   �      &           s_valid => _validW ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�+   �   �   �   �      %           s_valid => validW ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�/     �   �   �   �      '           m_ready => m_readyW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�/     �   �   �   �      &           m_ready => _readyW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�2   �   �   �   �      %           m_ready => readyW ( j+1 ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�7     �   �   �   �      '           s_ready => m_readyW ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�8     �   �   �   �      &           s_ready => _readyW ( j   ),5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^�9   �   �   �   �      %           s_ready => readyW ( j   ),5�_�  �  �  �      �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^��     �   y   �   �      u                  --if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo   B                  --   m_axis_tdata  <= wirex(ITER-1)(7 downto 0);   _                  --   m_axis_tvalid <= '1';                           --y ya no tengo mas nada   6                  --   state         <= waitingMready;   *                  --   bitCounter    := 0;                     --end if;5�_�  �  �          �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^��     �   y   {   �      s                  if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^��     �   y   {   �      r                  if _readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �  �      �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   y   {   �      q                  if readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   y       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�   �   x   y          Z                  m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   S       ����                                                                                                                                                                >   
                                                       �                                                                                              y          ~                 ^�5   �   R   S          !            readyW(0)     <= '1';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x          }                 ^�B   �   w   y   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              x          x          v       ^�H   �   w   y   �      q                  if readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   w       ����                                                                                                                                                                >   
                                                       �                                                                                              x          x          v       ^�3     �   v   x   �    �   w   x   �    5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�4     �   w   y   �      '                  validW(0)     <= '0';5�_�  �  �          �   x       ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�8     �   w   y   �      '                  readyW(0)     <= '0';5�_�  �  �          �   x   '    ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�Q     �   w   y   �      *                  readyW(ITER)     <= '0';5�_�  �  �          �   y       ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�     �   x   z   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   y       ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�3     �   x   z   �      n                  if validW(0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   y        ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�4    �   x   z   �      r                  if validW(ITER0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   z        ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�B     �   y   {   �    �   z   {   �    5�_�  �  �          �   z   '    ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�C     �   y   {   �      *                  readyW(ITER)     <= '1';5�_�  �  �          �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              y          y          v       ^�F     �   y   {          *                  readyW(ITER)     <= '0';5�_�  �  �          �   z        ����                                                                                                                                                                >   
                                                       �                                                                                              z          ~          V       ^�H  ! �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                        end if;�   �   �   �                           end case;�   �   �   �      &                        when others =>�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      "                           end if;�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                                 else�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      !                        when 2 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 1 =>�   �   �   �      '                     case bitCounter is�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      $               when waitingMready =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     state         <= waitingMready;�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   y   {   �      *                     readyW(ITER)  <= '0';�   x   z   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   w   y   �      *                  readyW(ITER)     <= '1';�   v   x   �      '                  validW(0)     <= '0';�   u   w   �      $               when waitingCordic =>�   t   v   �                        end if;�   s   u   �      2                     bitCounter := bitCounter + 1;�   r   t   �                           end case;�   q   s   �      &                        when others =>�   p   r   �      9                          state         <= waitingCordic;�   o   q   �      b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada�   n   p   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   m   o   �      /                          validW(0)     <= '1';�   l   n   �      !                          end if;�   k   m   �      :                                wirez(0) <= (others=>'0');�   j   l   �                                else �   i   k   �      $                             end if;�   h   j   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   g   i   �      "                             else �   f   h   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   e   g   �      8                             if s_axis_tdata(7)='1' then�   d   f   �      ,                          if inv(0)='1' then�   c   e   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   b   d   �      4                          wirey(0) <= (others=>'0');�   a   c   �      !                        when 1 =>�   `   b   �      !                          end if;�   _   a   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      5                          if s_axis_tdata(7)='1' then�   Y   [   �      4                          wirex(0) <= (others=>'0');�   X   Z   �      !                        when 0 =>�   W   Y   �      '                     case bitCounter is�   V   X   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   U   W   �      $               when waitingSvalid =>�   T   V   �                  case state is�   S   U   �               else�   R   T   �                  bitCounter    := 0;�   Q   S   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   P   R   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada�   O   Q   �      -            angle         <= (others => '0');�   N   P   �      !            clockWise     <= '0';�   M   O   �      -            m_axis_tdata  <= (others => '0');�   L   N   �      !            m_axis_tvalid <= '0';�   K   M   �      !            s_axis_tready <= '1';�   J   L   �      +            state         <= waitingSvalid;�   I   K   �               if rst = '0' then�   H   J   �            if rising_edge(clk) then�   G   I   �         begin�   F   H   �      9      variable extension :std_logic_vector (15 downto 0);�   E   G   �      *      variable sign :signed (15 downto 0);�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      %   cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      '   signal clockWise : std_logic := '0';�   5   7   �      "   signal xyData    : xyDataArray;�   4   6   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   y   {          -                     readyW(ITER)     <= '0';�   }             (                     bitCounter    := 0;�   |   ~          4                     state         <= waitingMready;�   {   }          ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   z   |          @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);5�_�  �  �          �   G       ����                                                                                                                                                                >   
                                                       �                                                                                                                               ^��     �   F   G          9      variable extension :std_logic_vector (15 downto 0);5�_�  �  �          �   E        ����                                                                                                                                                                >   
                                                       �                                                                                                                               ^��  " �   D   E           5�_�  �  �          �   C       ����                                                                                                                                                                >   
                                                       �                                                                                                                               ^��     �   B   D   �      %   cordic_proc:process (clk) is --{{{5�_�  �  �          �   C        ����                                                                                                                                                                >   
                                                       �                                                                                              C          �          V       ^��     �   B   �   �    �   C   D   �    5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �        !   end process cordic_proc; --}}}5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �        !   end process cordic_proc; --}}}5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �      5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �  	      )   pre_cordic_proc:process (clk) is --{{{5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �  	      %   end process pre_cordic_proc; --}}}5�_�  �  �          �   n       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�2     �   m   n          b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   W       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�`     �   V   X        !                        when 0 =>5�_�  �  �          �   `       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�c     �   _   a        !                        when 1 =>5�_�  �  �          �   q        ����                                                                                                                                                                >   
                                                       �                                                                                              q          q          V       ^�f     �   p   q          2                     bitCounter := bitCounter + 1;5�_�  �  �          �   V       ����                                                                                                                                                                >   
                                                       �                                                                                              q          q          V       ^�i     �   U   W      �   V   W      5�_�  �  �          �   v       ����                                                                                                                                                                >   
                                                       �                                                                                              r          r          V       ^��     �   u   w        q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   v       ����                                                                                                                                                                >   
                                                       �                                                                                              r          r          V       ^��     �   u   w        q                  if readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   v   !    ����                                                                                                                                                                >   
                                                       �                                                                                              r          r          V       ^��     �   v   x      5�_�  �  �          �   t        ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   s   t          '                  validW(0)     <= '0';5�_�  �  �          �   v        ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   u   w      �   v   w      5�_�  �  �          �   v       ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   u   w          '                  validW(0)     <= '0';5�_�  �  �          �   w        ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   v   x  	    �   w   x  	    5�_�  �  �          �   w       ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   v   x          k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo5�_�  �  �          �   w   '    ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   v   x  
      f                     s_axis_tready <= '0';                           --entonces yo tambien estoy listo5�_�  �  �          �   t       ����                                                                                                                                                                >   
                                                       �                                                                                              t          t          V       ^��     �   s   t          *                  readyW(ITER)     <= '1';5�_�  �  �          �   {        ����                                                                                                                                                                >   
                                                       �                                                                                              {          {          V       ^�     �   z   {          4                     state         <= waitingMready;5�_�  �  �          �   w        ����                                                                                                                                                                >   
                                                       �                                                                                              {          {          V       ^�     �   v   x      �   w   x      5�_�  �  �          �   w   -    ����                                                                                                                                                                >   
                                                       �                                                                                              |          |          V       ^�     �   v   x  	      4                     state         <= waitingMready;5�_�  �  �          �   |        ����                                                                                                                                                                >   
                                                       �                                                                                              |   '       |   '       V   2    ^�,     �   {   |          (                     bitCounter    := 0;5�_�  �  �          �   x        ����                                                                                                                                                                >   
                                                       �                                                                                              |   '       |   '       V   2    ^�-     �   w   y      �   x   y      5�_�  �  �  �      �   y        ����                                                                                                                                                                >   
                                                       �                                                                                              y           |           V        ^�V     �   x   y              *                     readyW(ITER)  <= '0';   @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);   ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada5�_�  �  �          �   z        ����                                                                                                                                                                >   
                                                       �                                                                                              z           �          V       ^�r     �   y   z              $               when waitingMready =>   l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   N                    bitCounter := bitCounter+1;                   --incremento   '                     case bitCounter is   !                        when 1 =>   E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);   !                        when 2 =>   3                           if(inv(ITER-1)='1') then   P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));   d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));                              else   O                              angle <= std_logic_vector(signed(wirez(ITER-1)));   I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);   "                           end if;   �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   0                           s_axis_tready <= '1';   .                           bitCounter    := 0;   �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato   &                        when others =>                        end case;5�_�  �  �          �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z           z          V       ^�s     �   y   z                            end if;5�_�  �  �          �   O   !    ����                                                                                                                                                                >   
                                                       �                                                                                              z           z          V       ^��     �   N   P   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   P   !    ����                                                                                                                                                                >   
                                                       �                                                                                              z           z          V       ^��     �   O   Q   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada5�_�  �  �          �   N       ����                                                                                                                                                                >   
                                                       �                                                                                              z           z          V       ^��     �   M   N          -            angle         <= (others => '0');5�_�  �  �          �   7       ����                                                                                                                                                                >   
                                                       �                                                                                              y           y          V       ^��     �   6   7          '   signal clockWise : std_logic := '0';5�_�  �  �          �   L       ����                                                                                                                                                                =   
                                                       �                                                                                              x           x          V       ^��     �   K   L          !            clockWise     <= '0';5�_�  �  �          �   �       ����                                                                                                                                                                =   
                                                       �                                                                                              w           w          V       ^��     �   �   �          !            clockWise     <= '0';5�_�  �  �          �   h        ����                                                                                                                                                                =   
                                                       �                                                                                              w           w          V       ^��     �   g   i          :                                wirez(0) <= (others=>'0');5�_�  �  �          �   K       ����                                                                                                                                                                =   
                                                       �                                                                                              w           w          V       ^��     �   J   K          -            m_axis_tdata  <= (others => '0');5�_�  �  �          �   J       ����                                                                                                                                                                =   
                                                       �                                                                                              v           v          V       ^��  # �   I   J          !            m_axis_tvalid <= '0';5�_�  �  �          �   4       ����                                                                                                                                                                =   
                                                       �                                                                                              u           u          V       ^��     �   3   5   �    �   4   5   �    5�_�  �             �   5   
    ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^��     �   4   6   �      1   signal state     : axiStates := waitingSvalid;5�_�  �                5       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^��     �   4   6   �      5   signal posSstate     : axiStates := waitingSvalid;5�_�                  5       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^��     �   4   6   �      4   signal posState     : axiStates := waitingSvalid;5�_�                 5       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^��     �   4   6   �      3   signal posState    : axiStates := waitingSvalid;5�_�                 5       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^�      �   4   6   �      2   signal posState   : axiStates := waitingSvalid;5�_�                 }       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^�     �   |   }          *      variable sign :signed (15 downto 0);5�_�                 E       ����                                                                                                                                                                >   
                                                       �                                                                                              v           v          V       ^�     �   D   E          *      variable sign :signed (15 downto 0);5�_�                        ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�#     �   ~   �   �      +            state         <= waitingSvalid;5�_�                        ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�&     �   ~   �   �      /            posSstate         <= waitingSvalid;5�_�    	                    ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�(     �   ~   �   �      .            posState         <= waitingSvalid;5�_�    
          	   �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�.     �      �          !            s_axis_tready <= '1';5�_�  	            
   �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�J     �   �   �   �      T            validW(0)     <= '0';                           --y ya no tengo mas nada5�_�  
               �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�[     �   �   �   �      T            readyW(0)     <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�`     �   �   �   �      W            readyW(ITER)     <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�`     �   �   �   �      V            readyW(ITER)    <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�`     �   �   �   �      U            readyW(ITER)   <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^�l     �   �   �   �      T            readyW(ITER)  <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^��     �   �   �          T            inv(0)        <= '0';                           --y ya no tengo mas nada5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^��     �   �   �   �                  bitCounter    := 0;5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              u           u          V       ^��     �   �   �   �      #            posBbitCounter    := 0;5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �          '                     case bitCounter is5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �          !                        when 0 =>5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      5                          if s_axis_tdata(7)='1' then5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      4                          f s_axis_tdata(7)='1' then5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      3                           s_axis_tdata(7)='1' then5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      2                          s_axis_tdata(7)='1' then5�_�                 �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^��     �   �   �   �      2                          m_axis_tdata(7)='1' then5�_�                 �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^�     �   �   �   �      2                          m_axis_tdata(7)='1' then5�_�                 �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^�     �   �   �   �      1                          m_axis_tdata7)='1' then5�_�                 �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^�     �   �   �   �      0                          m_axis_tdata)='1' then5�_�                 �   '    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �   !       v   !    ^�     �   �   �   �      /                          m_axis_tdata='1' then5�_�                  �        ����                                                                                                                                                                >   
                                                       �                                                                                              �           �           V        ^�l     �   �   �   �    �   �   �   �    �   �   �          '                          m_axis_tdata=5�_�    !              �        ����                                                                                                                                                                >   
                                                       �                                                                                              �           �           V        ^��     �   �   �   �    �   �   �   �    �   �   �          P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));   d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));                              else   O                              angle <= std_logic_vector(signed(wirez(ITER-1)));   I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);5�_�     "          !   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          4                          wirex(0) <= (others=>'0');5�_�  !  #          "   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          -                             inv(0)   <= '1';5�_�  "  $          #   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));5�_�  #  %          $   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �                                    else5�_�  $  &          %   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          -                             inv(0)   <= '0';5�_�  %  '          &   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));5�_�  &  (          '   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   !       V        ^��     �   �   �          !                          end if;5�_�  '  )          (   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          "                           end if;�   �   �          I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �          O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �                                     else�   �   �          d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �          P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �          3                           if(inv(ITER-1)='1') then5�_�  (  *          )   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �    5�_�  )  +          *   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �                           �   �   �   �    5�_�  *  ,          +   �   (    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �    �   �   �   �    5�_�  +  -          ,   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�H     �   �   �   �      )                     m_axis_tvalid = '1';5�_�  ,  .          -   �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�J     �   �   �   �      )                     m_axis_tready = '1';5�_�  -  /          .   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�\     �   �   �   �    �   �   �   �    5�_�  .  0          /   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�]     �   �   �          "            posBitCounter    := 0;5�_�  /  1          0   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�^     �   �   �   �                           �   �   �   �    5�_�  0  2          1   �   .    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�t     �   �   �   �                           �   �   �   �    5�_�  1  3          2   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �           V       ^��     �   �   �          !                        when 1 =>   4                          wirey(0) <= (others=>'0');   g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));   ,                          if inv(0)='1' then   8                             if s_axis_tdata(7)='1' then   _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));   "                             else    `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));   $                             end if;                             else    :                                wirez(0) <= (others=>'0');   !                          end if;   /                          validW(0)     <= '1';   k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo   b                          m_axis_tvalid <= '0';                           --y ya no tengo mas nada   9                          state         <= waitingCordic;   &                        when others =>                        end case;   2                     bitCounter := bitCounter + 1;                     end if;   $               when waitingCordic =>   '                  validW(0)     <= '0';   *                  readyW(ITER)     <= '1';   q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo   *                     readyW(ITER)  <= '0';   @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);   ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada   4                     state         <= waitingMready;   (                     bitCounter    := 0;                     end if;    5�_�  2  4          3   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          $               when waitingMready =>   l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   N                    bitCounter := bitCounter+1;                   --incremento   '                     case bitCounter is   !                        when 1 =>   E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);   !                        when 2 =>   3                           if(inv(ITER-1)='1') then   P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));   d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));                              else   O                              angle <= std_logic_vector(signed(wirez(ITER-1)));   I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);   "                           end if;5�_�  3  5          4   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �    �   �   �   �    5�_�  4  6          5   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �                           �   �   �   �    5�_�  5  7          6   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �           5�_�  6  8          7   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �           5�_�  7  9          8   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �           5�_�  8  :          9   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          .                           bitCounter    := 0;5�_�  9  ;          :   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  :  <          ;   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �                                 �   �   �   �    5�_�  ;  =          <   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          &                        when others =>5�_�  <  >          =   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �                               end case;5�_�  =  ?          >   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �                            end if;5�_�  >  @          ?   �   
    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �                      end case;5�_�  ?  A          @   �   	    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �                   end if;5�_�  @  B          A   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �                end if;5�_�  A  C          B           ����                                                                                                                                                                >   
                                                       �                                                                                                 	       �   	       V   	    ^��     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                              end if;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �      /                     posState := waitingMready;�   �   �   �      +                     posBitCounter    := 0;�   �   �   �      )                     m_axis_tready = '0';�   �   �   �      )                     m_axis_tvalid = '1';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case state is�   �   �   �               else�   �   �   �                  posBitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�      �   �      !            m_axis_tvalid <= '0';�   ~   �   �      +            posState      <= waitingSvalid;�   }      �               if rst = '0' then�   |   ~   �            if rising_edge(clk) then�   {   }   �         begin�   z   |   �      1      variable bitCounter :integer range 0 to 8 ;�   y   {   �      )   pos_cordic_proc:process (clk) is --{{{�   w   y   �      %   end process pre_cordic_proc; --}}}�   v   x   �            end if;�   u   w   �               end if;�   t   v   �                  end case;�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     state         <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingCordic =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          state         <= waitingCordic;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case state is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            state         <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   ~   �          +            posState      <= waitingSvalid;�   �   �          "            posBitCounter    := 0;�   �   �          -            m_axis_tdata  <= (others => '0');�      �          !            m_axis_tvalid <= '0';�   �   �          T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �          -            angle         <= (others => '0');5�_�  B  D          C   �       ����                                                                                                                                                                >   
                                                       �                                                                                                 	       �   	       V   	    ^�     �   �   �   �                  case state is5�_�  C  E          D   �       ����                                                                                                                                                                >   
                                                       �                                                                                                 	       �   	       V   	    ^�     �   �   �   �                  case posSstate is5�_�  D  F          E   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                              end if;�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �      4                     posState      := waitingMready;�   �   �   �      (                     posBitCounter := 0;�   �   �   �      *                     m_axis_tready  = '0';�   �   �   �      *                     m_axis_tvalid  = '1';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  posBitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�      �   �      !            m_axis_tvalid <= '0';�   ~   �   �      +            posState      <= waitingSvalid;�   }      �               if rst = '0' then�   |   ~   �            if rising_edge(clk) then�   {   }   �         begin�   z   |   �      1      variable bitCounter :integer range 0 to 8 ;�   y   {   �      )   pos_cordic_proc:process (clk) is --{{{�   w   y   �      %   end process pre_cordic_proc; --}}}�   v   x   �            end if;�   u   w   �               end if;�   t   v   �                  end case;�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     state         <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingCordic =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          state         <= waitingCordic;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case state is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            state         <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          )                     m_axis_tvalid = '1';�   �   �          /                     posState := waitingMready;�   �   �          +                     posBitCounter    := 0;�   �   �          )                     m_axis_tready = '0';5�_�  E  G          F   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�#     �   �   �          0                           s_axis_tready <= '1';�   �   �          �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �          �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �          .                           bitCounter    := 0;5�_�  F  H          G   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�%     �   �   �                                  end if;5�_�  G  J          H   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�/     �   �   �   �      -                        s_axis_tready <= '1';5�_�  H  L  I      J   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�e     �   �   �   �                           �   �   �   �    5�_�  J  M  K      L   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �          *                     m_axis_tready  = '0';5�_�  L  N          M   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �    �   �   �   �    �   �   �          -                        m_axis_tready <= '1';5�_�  M  O          N   �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   (       V       ^��     �   �   �   �      )                     readyW(ITER) := '0';5�_�  N  P          O   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �           �   (       V       ^��     �   �   �          )                     readyW(ITER) := '1';5�_�  O  Q          P   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  := '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �      4                     posState      := waitingMready;�   �   �   �      (                     posBitCounter := 0;�   �   �   �      *                     m_axis_tvalid  = '1';�   �   �   �      )                     readyW(ITER) := '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  posBitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�      �   �      !            m_axis_tvalid <= '0';�   ~   �   �      +            posState      <= waitingSvalid;�   }      �               if rst = '0' then�   |   ~   �            if rising_edge(clk) then�   {   }   �         begin�   z   |   �      1      variable bitCounter :integer range 0 to 8 ;�   y   {   �      )   pos_cordic_proc:process (clk) is --{{{�   w   y   �      %   end process pre_cordic_proc; --}}}�   v   x   �            end if;�   u   w   �               end if;�   t   v   �                  end case;�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     state         <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingCordic =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          state         <= waitingCordic;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case state is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            state         <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          +                        bitCounter    := 0;�   �   �          ,                        readyW(ITER) := '1';�   �   �          �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �          }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  P  R          Q   �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  := '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �      4                     posState      := waitingMready;�   �   �   �      (                     posBitCounter := 0;�   �   �   �      *                     m_axis_tvalid  = '1';�   �   �   �      *                     readyW(ITER)  := '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  posBitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�      �   �      !            m_axis_tvalid <= '0';�   ~   �   �      +            posState      <= waitingSvalid;�   }      �               if rst = '0' then�   |   ~   �            if rising_edge(clk) then�   {   }   �         begin�   z   |   �      1      variable bitCounter :integer range 0 to 8 ;�   y   {   �      )   pos_cordic_proc:process (clk) is --{{{�   w   y   �      %   end process pre_cordic_proc; --}}}�   v   x   �            end if;�   u   w   �               end if;�   t   v   �                  end case;�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     state         <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingCordic =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          state         <= waitingCordic;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case state is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            state         <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal state     : axiStates := waitingSvalid;�   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          )                     readyW(ITER) := '0';�   �   �          4                     posState      := waitingMready;�   �   �          (                     posBitCounter := 0;�   �   �          *                     m_axis_tvalid  = '1';5�_�  Q  S          R   �   #    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �      *                     m_axis_tvalid  = '1';5�_�  R  T          S   4   
    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   3   5   �      1   signal state     : axiStates := waitingSvalid;5�_�  S  U          T   4       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   3   5   �      5   signal preSstate     : axiStates := waitingSvalid;5�_�  T  V          U   4       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   3   5   �      4   signal preState     : axiStates := waitingSvalid;5�_�  U  W          V   4       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   3   5   �      3   signal preState    : axiStates := waitingSvalid;5�_�  V  Z          W   4       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�   $ �   3   5   �      2   signal preState   : axiStates := waitingSvalid;5�_�  W  [  X      Z   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  Z  \          [   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�  % �   �   �                               end if;5�_�  [  ]          \   H       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�     �   G   I   �      +            state         <= waitingSvalid;5�_�  \  ^          ]   H       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�      �   G   I   �      /            preSstate         <= waitingSvalid;5�_�  ]  _          ^   H       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�"     �   G   I   �      .            preState         <= waitingSvalid;5�_�  ^  `          _   H       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�#  & �   G   I   �      *            preState     <= waitingSvalid;5�_�  _  a          `   N       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�'     �   M   O   �                  case state is5�_�  `  b          a   N       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�)  ( �   M   O   �                  case preSstate is5�_�  a  c          b   k       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�^     �   j   l   �    �   k   l   �    5�_�  b  d          c   k       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�`  ) �   j   l   �      &                        when others =>5�_�  c  e          d   k        ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�m     �   j   k          -                        when waitingMready =>5�_�  d  f          e   u       ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�r     �   t   v   �    �   u   v   �    5�_�  e  g          f   u       ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�s  * �   t   v          &                        when others =>5�_�  f  h          g   j       ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�x     �   i   k   �      9                          state         <= waitingCordic;5�_�  g  i          h   j       ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�z     �   i   k   �      =                          preSstate         <= waitingCordic;5�_�  h  j          i   j   (    ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^�{  + �   i   k   �      <                          preState         <= waitingCordic;5�_�  i  k          j   j   2    ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^��     �   i   k   �      9                          preState      <= waitingCordic;5�_�  j  l          k   n       ����                                                                                                                                                                >   
                                                       �                                                                                              k          k          V       ^��     �   m   o   �      $               when waitingCordic =>5�_�  k  m          l   3   6    ����                                                                                                                                                                >   
                                                       �                                                                                              3   6       3   C       v   C    ^��  , �   2   4   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);5�_�  l  n          m   r       ����                                                                                                                                                                >   
                                                       �                                                                                              3   6       3   C       v   C    ^��     �   q   s   �      4                     state         <= waitingSvalid;5�_�  m  o          n   r       ����                                                                                                                                                                >   
                                                       �                                                                                              3   6       3   C       v   C    ^��     �   q   s   �      8                     preSstate         <= waitingSvalid;5�_�  n  p          o   p        ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�  - �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  := '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      := waitingMready;�   �   �   �      (                     posBitCounter := 0;�   �   �   �      *                     m_axis_tvalid := '1';�   �   �   �      *                     readyW(ITER)  := '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  posBitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�      �   �      +            posState      <= waitingSvalid;�   ~   �   �               if rst = '0' then�   }      �            if rising_edge(clk) then�   |   ~   �         begin�   {   }   �      1      variable bitCounter :integer range 0 to 8 ;�   z   |   �      )   pos_cordic_proc:process (clk) is --{{{�   x   z   �      %   end process pre_cordic_proc; --}}}�   w   y   �            end if;�   v   x   �               end if;�   u   w   �                  end case;�   t   v   �                     when others =>�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     preState      <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingMready =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          preState      <= waitingMready;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case preState is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            preState      <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   o   q          *                     validW(0)     <= '0';�   r   t          (                     bitCounter    := 0;�   q   s          7                     preState         <= waitingSvalid;�   p   r          f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo5�_�  o  q          p   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�     �   �   �   �                  posBitCounter := 0;5�_�  p  r          q   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�     �   �   �   �                  osBitCounter := 0;5�_�  q  s          r   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�     �   �   �   �                  sBitCounter := 0;5�_�  r  t          s   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�  . �   �   �   �                  BitCounter := 0;5�_�  s  u          t   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�)     �   �   �   �      *                     readyW(ITER)  := '0';5�_�  t  v          u   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�*  / �   �   �   �      )                     ready(ITER)  := '0';5�_�  u  w          v   >       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�P     �   =   ?   �      A   signal validW,  readyW,inv  : handShakeVector:= (others=>'0');5�_�  v  x          w   >       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�Q  0 �   =   ?   �      @   signal validW, readyW,inv  : handShakeVector:= (others=>'0');5�_�  w  y          x   >       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^�Y  3 �   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');5�_�  x  z          y   �   #    ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��  4 �   �   �   �      *                     readyW(ITER)  := '0';5�_�  y  {          z   �   #    ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��  5 �   �   �   �      *                     m_axis_tvalid := '1';5�_�  z  |          {   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��     �   �   �   �      (                     posBitCounter := 0;5�_�  {  }          |   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��     �   �   �   �      '                     osBitCounter := 0;5�_�  |  ~          }   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��     �   �   �   �      &                     sBitCounter := 0;5�_�  }            ~   �       ����                                                                                                                                                                >   
                                                       �                                                                                              p           s           V        ^��  6 �   �   �   �      %                     BitCounter := 0;5�_�  ~  �             �        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��  7 �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  := '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      := waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�      �   �      +            posState      <= waitingSvalid;�   ~   �   �               if rst = '0' then�   }      �            if rising_edge(clk) then�   |   ~   �         begin�   {   }   �      1      variable bitCounter :integer range 0 to 8 ;�   z   |   �      )   pos_cordic_proc:process (clk) is --{{{�   x   z   �      %   end process pre_cordic_proc; --}}}�   w   y   �            end if;�   v   x   �               end if;�   u   w   �                  end case;�   t   v   �                     when others =>�   s   u   �                        end if;�   r   t   �      (                     bitCounter    := 0;�   q   s   �      4                     preState      <= waitingSvalid;�   p   r   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   o   q   �      *                     validW(0)     <= '0';�   n   p   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   m   o   �      $               when waitingMready =>�   l   n   �                        end if;�   k   m   �                           end case;�   j   l   �      &                        when others =>�   i   k   �      9                          preState      <= waitingMready;�   h   j   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   g   i   �      /                          validW(0)     <= '1';�   f   h   �      !                          end if;�   e   g   �      7                             wirez(0) <= (others=>'0');�   d   f   �                                else �   c   e   �      $                             end if;�   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   a   c   �      "                             else �   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   _   a   �      8                             if s_axis_tdata(7)='1' then�   ^   `   �      ,                          if inv(0)='1' then�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   \   ^   �      4                          wirey(0) <= (others=>'0');�   [   ]   �      !                        when 2 =>�   Z   \   �      !                          end if;�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   X   Z   �      -                             inv(0)   <= '0';�   W   Y   �                                else�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   U   W   �      -                             inv(0)   <= '1';�   T   V   �      5                          if s_axis_tdata(7)='1' then�   S   U   �      4                          wirex(0) <= (others=>'0');�   R   T   �      !                        when 1 =>�   Q   S   �      '                     case bitCounter is�   P   R   �      2                     bitCounter := bitCounter + 1;�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   N   P   �      $               when waitingSvalid =>�   M   O   �                  case preState is�   L   N   �               else�   K   M   �                  bitCounter    := 0;�   J   L   �      !            inv(0)        <= '0';�   I   K   �      !            validW(0)     <= '0';�   H   J   �      !            s_axis_tready <= '1';�   G   I   �      +            preState      <= waitingSvalid;�   F   H   �               if rst = '0' then�   E   G   �            if rising_edge(clk) then�   D   F   �         begin�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          *                     readyW(ITER)  <= '0';�   �   �          4                     posState      := waitingMready;�   �   �          %                     bitCounter := 0;�   �   �          *                     m_axis_tvalid <= '1';5�_�    �          �   �   #    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��  8 �   �   �   �      4                     posState      := waitingMready;5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �      }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  �  �          �   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �      �                        posSstate         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  �  �          �   �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��  9 �   �   �   �      �                        posState         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  �  �          �   �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �   �      -                        readyW(ITER)  := '1';5�_�  �  �          �   �   &    ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��  < �   �   �   �      -                        readyW(ITER)  M= '1';5�_�  �  �  �      �   @       ����                                                                                                                                                                >   
                                                       �                                                                                                                               ^�     �   ?   A   �    �   @   A   �    5�_�  �  �          �   A       ����                                                                                                                                                                >   
                                                       �                                                                                                                               ^�     �   @   A          j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   >        ����                                                                                                                                                                >   
                                                       �                                                                                              >          >          V       ^�)     �   =   >          A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');5�_�  �  �          �   <       ����                                                                                                                                                                    
                                                       �                                                                                              >          >          V       ^�*     �   ;   =   �    �   <   =   �    5�_�  �  �          �   :        ����                                                                                                                                                                    
                                                       �                                                                                              ?          ?          V       ^�-     �   9   =   �       5�_�  �  �          �   <        ����                                                                                                                                                                    
                                                       �                                                                                              A          A          V       ^     �   ;   <           5�_�  �  �          �   =       ����                                                                                                                                                                    
                                                       �                                                                                              @          @          V       ^     �   =   ?   �    5�_�  �  �          �   @       ����                                                                                                                                                                    
                                                       �                                                                                              A          A          V       ^     �   ?   A   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   @   #    ����                                                                                                                                                                    
                                                       �                                                                                              A          A          V       ^     �   ?   A   �      �   type   intLUT        is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   ?   4    ����                                                                                                                                                                    
                                                       �                                                                                              A          A          V       ^     �   >   @   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);5�_�  �  �          �   @   E    ����                                                                                                                                                                    
                                                       �                                                                                              A          A          V       ^     �   ?   A   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   ?   M    ����                                                                                                                                                                    
                                                       �                                                                                              @   M       ?   M          M    ^¤     �   ?   A   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer         range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   >   @   �      \   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector(N-1 downto 0);5�_�  �  �          �   A       ����                                                                                                                                                                    
                                                       �                                                                                              @   M       ?   M          M    ^­     �   A   C   �    5�_�  �  �          �   >        ����                                                                                                                                                                    
                                                       �                                                                                              @   M       ?   M          M    ^¯     �   =   @   �       5�_�  �  �          �   A        ����                                                                                                                                                                    
                                                       �                                                                                              A   (       A   (       V   (    ^��     �   @   A          �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   C       ����                                                                                                                                                                    
                                                       �                                                                                              A   (       A   (       V   (    ^��     �   B   D   �    �   C   D   �    5�_�  �  �          �   ?       ����                                                                                                                                                                    
                                                       �                                                                                              A   (       A   (       V   (    ^��     �   >   @   �      	   --con 5�_�  �  �          �   ?       ����                                                                                                                                                                    
                                                       �                                                                                              A   (       A   (       V   (    ^��     �   >   @   �         --5�_�  �  �          �   ?   
    ����                                                                                                                                                                    
                                                       �                                                                                              A   (       A   (       V   (    ^��     �   ?   A   �         �   ?   A   �    5�_�  �  �          �   D   7    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   C   E   �         �   C   E   �    5�_�  �  �          �   D   G    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�     �   C   E   �      G   --defino una tabla con los angulos tal que su arcotangente da 1/2**N5�_�  �  �          �   V   .    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�q     �   U   W   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   V   .    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�r     �   U   W   �      .                  if s_axis_tvalid = '1' then 5�_�  �  �          �   W   2    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�~     �   V   X   �      2                     bitCounter := bitCounter + 1;5�_�  �  �          �   [   5    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   Z   \   �      5                          if s_axis_tdata(7)='1' then5�_�  �  �          �   [   6    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   Z   \   �      6                          if s_axis_tdata(7)='1' then 5�_�  �  �          �   ]   f    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   \   ^   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));5�_�  �  �          �   `   e    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   _   a   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));5�_�  �  �          �   d   b    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   c   e   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));5�_�  �  �          �   Z       ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   Y   Z          4                          wirex(0) <= (others=>'0');5�_�  �  �          �   Z   ;    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   Y   [   �      B                          if s_axis_tdata(7)='1' then    --si el x5�_�  �  �          �   Z   ;    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   Y   [   �      ;                          if s_axis_tdata(7)='1' then    --5�_�  �  �          �   Y   !    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�     �   X   Z   �      !                        when 1 =>5�_�  �  �          �   Y   "    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�     �   X   Z   �      $                        when 1 => --5�_�  �  �          �   Y   ;    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�     �   X   Z   �      ;                        when 1 =>                        --5�_�  �  �          �   b       ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��     �   a   b          4                          wirey(0) <= (others=>'0');5�_�  �  �          �   a   !    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^��  = �   `   b   �      !                        when 2 =>5�_�  �  �          �   c   ,    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�     �   b   d   �      ,                          if inv(0)='1' then5�_�  �  �          �   m   5    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�V     �   m   p   �                                �   m   o   �    5�_�  �  �          �   n   (    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�j     �   m   o   �      )                          if readyW(0) = 5�_�  �  �          �   o       ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�r     �   n   o                                    15�_�  �  �          �   a   "    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�Q     �   `   b   �      :                        when 2 => --el y se copia tal cual5�_�  �  �          �   c   -    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^�Y     �   b   d   �      z                          if inv(0)='1' then --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z5�_�  �  �          �   n   +    ����                                                                                                                                                                    
                                                       �                                                                                              B   (       B   (       V   (    ^Ӛ     �   m   o   �      -                          if readyW(0) ='1'  5�_�  �  �          �   V   9    ����                                                                                                                                                                    
                                                       �                                                                                              V   9       Z   9          9    ^��     �   V   [   �      g                     bitCounter := bitCounter + 1;       --espero 2 datos de 8 bits.. primero X luego Y   '                     case bitCounter is   <                        when 1 =>                        --X   q                          if s_axis_tdata(7)='1' then    --corrijo cuadrante si X es negativo y lo informo en inv�   U   W   �      T                  if s_axis_tvalid = '1' then            --espero a que entren datos5�_�  �  �          �   a   9    ����                                                                                                                                                                    
                                                       �                                                                                              V   9       Z   9          9    ^��     �   `   b   �      Q                        when 2 =>                        --el y se copia tal cual5�_�  �  �          �   c   9    ����                                                                                                                                                                    
                                                       �                                                                                              V   9       Z   9          9    ^��     �   b   d   �      �                          if inv(0)='1' then             --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z5�_�  �  �          �   m   J    ����                                                                                                                                                                    
                                                       �                                                                                              V   9       Z   9          9    ^�     �   l   n   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo5�_�  �  �          �   o       ����                                                                                                                                                                    
                                                       �                                                                                              V   9       Z   9          9    ^�5     �   n   p   �      9                          preState      <= waitingMready;5�_�  �  �          �   o        ����                                                                                                                                                                    
                                                       �                                                                                              o   )       o   )       V   )    ^�<     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�      �   �      )   pos_cordic_proc:process (clk) is --{{{�   }      �      %   end process pre_cordic_proc; --}}}�   |   ~   �            end if;�   {   }   �               end if;�   z   |   �                  end case;�   y   {   �                     when others =>�   x   z   �                        end if;�   w   y   �      (                     bitCounter    := 0;�   v   x   �      4                     preState      <= waitingSvalid;�   u   w   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   t   v   �      *                     validW(0)     <= '0';�   s   u   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   r   t   �      $               when waitingMready =>�   q   s   �                        end if;�   p   r   �                           end case;�   o   q   �      &                        when others =>�   n   p   �      =                              preState      <= waitingMready;�   m   o   �      +                          if readyW(0) ='1'�   l   n   �      �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo�   k   m   �      /                          validW(0)     <= '1';�   j   l   �      !                          end if;�   i   k   �      7                             wirez(0) <= (others=>'0');�   h   j   �                                else �   g   i   �      $                             end if;�   f   h   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   e   g   �      "                             else �   d   f   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   c   e   �      8                             if s_axis_tdata(7)='1' then�   b   d   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   a   c   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      �                        when 2 =>                                                                           --el y se copia tal cual�   _   a   �      !                          end if;�   ^   `   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '0';�   \   ^   �                                else�   [   ]   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   Z   \   �      -                             inv(0)   <= '1';�   Y   [   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   n   p          =                              preState      <= waitingMready;5�_�  �  �          �   o        ����                                                                                                                                                                    
                                                       �                                                                                              o           o           V        ^�>  > �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�      �   �      )   pos_cordic_proc:process (clk) is --{{{�   }      �      %   end process pre_cordic_proc; --}}}�   |   ~   �            end if;�   {   }   �               end if;�   z   |   �                  end case;�   y   {   �                     when others =>�   x   z   �                        end if;�   w   y   �      (                     bitCounter    := 0;�   v   x   �      4                     preState      <= waitingSvalid;�   u   w   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   t   v   �      *                     validW(0)     <= '0';�   s   u   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   r   t   �      $               when waitingMready =>�   q   s   �                        end if;�   p   r   �                           end case;�   o   q   �      &                        when others =>�   n   p   �      8                              preState <= waitingMready;�   m   o   �      +                          if readyW(0) ='1'�   l   n   �      �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo�   k   m   �      /                          validW(0)     <= '1';�   j   l   �      !                          end if;�   i   k   �      7                             wirez(0) <= (others=>'0');�   h   j   �                                else �   g   i   �      $                             end if;�   f   h   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   e   g   �      "                             else �   d   f   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   c   e   �      8                             if s_axis_tdata(7)='1' then�   b   d   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   a   c   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      �                        when 2 =>                                                                           --el y se copia tal cual�   _   a   �      !                          end if;�   ^   `   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '0';�   \   ^   �                                else�   [   ]   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   Z   \   �      -                             inv(0)   <= '1';�   Y   [   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   n   p          =                              preState      <= waitingMready;5�_�  �  �          �   v   D    ����                                                                                                                                                                    
                                                       �                                                                                              o           o           V        ^Ԯ  ? �   u   w   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo5�_�  �  �          �   n   +    ����                                                                                                                                                                    
                                                       �                                                                                              v   D       u   *          D    ^Զ  @ �   m   o   �      +                          if readyW(0) ='1'5�_�  �  �          �   p       ����                                                                                                                                                                    
                                                       �                                                                                              v   D       u   *          D    ^��  B �   o   q   �    �   p   q   �    5�_�  �  �          �   F       ����                                                                                                                                                                    
                                                       �                                                                                              w   D       v   *          D    ^�9  C �   E   G   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   l   /    ����                                                                                                                                                                    
                                                       �                                                                                              w   D       v   *          D    ^�P     �   k   m   �      /                          validW(0)     <= '1';5�_�  �  �          �   l   0    ����                                                                                                                                                                    
                                                       �                                                                                              w   D       v   *          D    ^�]     �   k   m   �      j                          validW(0)     <= '1'; --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   p        ����                                                                                                                                                                    
                                                       �                                                                                              v   &       y   &       V   &    ^�h     �   o   t   �    �   p   q   �    5�_�  �  �          �   p        ����                                                                                                                                                                    
                                                       �                                                                                              p          s          V       ^�k     �   r   t          (                     bitCounter    := 0;�   q   s          4                     preState      <= waitingSvalid;�   p   r          e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   o   q          *                     validW(0)     <= '0';5�_�  �  �          �   Z   *    ����                                                                                                                                                                    
                                                       �                                                                                              p          s          V       ^ռ     �   Y   [   �    �   Z   [   �    5�_�  �  �          �   Z   ,    ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^տ     �   Y   [   �      �                          validW(0)     <= '1';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   Z   ,    ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^��     �   Y   [   �      �                          validW(0)     <= '-';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   w       ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^��     �   w   z   �                           �   w   y   �    5�_�  �  �          �   y        ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^��     �   y   {   �    �   y   z   �    5�_�  �  �          �   y        ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^��     �   x   y           5�_�  �  �          �   y       ����                                                                                                                                                                    
                                                       �                                                                                              q          t          V       ^��     �   x   z          �                          validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   y        ����                                                                                                                                                                    
                                                       �                                                                                              y   $       y   $       V   $    ^��     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                     when others =>�   �   �   �                        end if;�      �   �      (                     bitCounter    := 0;�   ~   �   �      4                     preState      <= waitingSvalid;�   }      �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   |   ~   �      *                     validW(0)     <= '0';�   {   }   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   z   |   �      $               when waitingMready =>�   y   {   �                        end if;�   x   z   �      `                     validW(0) <= '0';--aviso al primero del pipeline que tengo los datos listos�   w   y   �                        else�   v   x   �                           end case;�   u   w   �      &                        when others =>�   t   v   �      !                          end if;�   s   u   �      1                              bitCounter    := 0;�   r   t   �      =                              preState      <= waitingSvalid;�   q   s   �      n                              s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   p   r   �      3                              validW(0)     <= '0';�   o   q   �      8                              preState <= waitingMready;�   n   p   �      0                          if readyW(0) ='1' then�   m   o   �      �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo�   l   n   �      �                          validW(0)     <= '1';                                                             --aviso al primero del pipeline que tengo los datos listos�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      �                          validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   x   z          �                     validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   y   &    ����                                                                                                                                                                    
                                                       �                                                                                              y   $       y   $       V   $    ^��     �   x   z   �      `                     validW(0) <= '0';--aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   s        ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^��     �   s   u   �    5�_�  �  �          �   u       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^��     �   u   w   �                                    �   u   w   �    5�_�  �  �          �   w       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^��     �   v   x   �    �   w   x   �    5�_�  �  �          �   t        ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�     �   s   t           5�_�  �  �          �   p       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�     �   o   p          8                              preState <= waitingMready;5�_�  �  �          �   p       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�     �   o   p          3                              validW(0)     <= '0';5�_�  �  �          �   q       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�+     �   p   q          =                              preState      <= waitingSvalid;5�_�  �  �          �   s       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�7     �   r   t   �    �   s   t   �    5�_�  �  �          �   s       ����                                                                                                                                                                    
                                                       �                                                                                              p   )       p   )       V   )    ^�:     �   r   t          �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo5�_�  �  �          �   s        ����                                                                                                                                                                    
                                                       �                                                                                              s          t          V       ^�>     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�   �   �   �                     when others =>�   �   �   �                        end if;�      �   �      (                     bitCounter    := 0;�   ~   �   �      4                     preState      <= waitingSvalid;�   }      �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   |   ~   �      *                     validW(0)     <= '0';�   {   }   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   z   |   �      $               when waitingMready =>�   y   {   �                        end if;�   x   z   �      &                     validW(0) <= '0';�   w   y   �                        else�   v   x   �                           end case;�   u   w   �      &                        when others =>�   t   v   �      !                          end if;�   s   u   �      =                              preState      <= waitingMready;�   r   t   �      T                              s_axis_tready <= '0';--entonces yo tambien estoy listo�   q   s   �                                  else �   p   r   �      1                              bitCounter    := 0;�   o   q   �      n                              s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   n   p   �      0                          if readyW(0) ='1' then�   m   o   �      �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo�   l   n   �      �                          validW(0)     <= '1';                                                             --aviso al primero del pipeline que tengo los datos listos�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      �                          validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   r   t          �                              s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo�   s   u          8                              preState <= waitingMready;5�_�  �  �          �   s   3    ����                                                                                                                                                                    
                                                       �                                                                                              s          t          V       ^�@     �   r   t   �      T                              s_axis_tready <= '0';--entonces yo tambien estoy listo5�_�  �  �          �   n       ����                                                                                                                                                                    
                                                       �                                                                                              s          t          V       ^�D     �   m   n          �                          s_axis_tready <= '0';                                                             --entonces yo tambien estoy listo5�_�  �  �          �   o       ����                                                                                                                                                                    
                                                       �                                                                                              r          s          V       ^�F     �   n   o          n                              s_axis_tready <= '1';                          --entonces yo tambien estoy listo5�_�  �  �          �   m        ����                                                                                                                                                                    
                                                       �                                                                                              m          m          V       ^�K     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      =                              preState      <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      1                              bitCounter    := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      e                          validW(0) <= '1';--aviso al primero del pipeline que tengo los datos listos�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      �                          validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   l   n          �                          validW(0)     <= '1';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   m   +    ����                                                                                                                                                                    
                                                       �                                                                                              m          m          V       ^�P     �   l   n   �      e                          validW(0) <= '1';--aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   Z        ����                                                                                                                                                                    
                                                       �                                                                                              Z   '       Z   '       V   '    ^�o     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      =                              preState      <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      1                              bitCounter    := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      +                          validW(0) <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      e                          validW(0) <= '0';--aviso al primero del pipeline que tengo los datos listos�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   Y   [          �                          validW(0)     <= '0';                                                             --aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   Z   +    ����                                                                                                                                                                    
                                                       �                                                                                              Z   '       Z   '       V   '    ^�r     �   Y   [   �      e                          validW(0) <= '0';--aviso al primero del pipeline que tengo los datos listos5�_�  �  �          �   r        ����                                                                                                                                                                    
                                                       �                                                                                              r   (       r   (       V   (    ^�~     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      8                              preState <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      1                              bitCounter    := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      +                          validW(0) <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      +                          validW(0) <= '0';�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   q   s          =                              preState      <= waitingMready;5�_�  �  �  �      �   q        ����                                                                                                                                                                    
                                                       �                                                                                              q          r          V       ^ւ  D �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      =                              preState      <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      1                              bitCounter    := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      +                          validW(0) <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      +                          validW(0) <= '0';�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   p   r          3                              s_axis_tready <= '0';�   q   s          8                              preState <= waitingMready;5�_�  �  �          �   o        ����                                                                                                                                                                    
                                                       �                                                                                              o          o          V       ^֢     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      =                              preState      <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      1                              bitCounter    := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      +                          validW(0) <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      +                          validW(0) <= '0';�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   n   p          1                              bitCounter    := 0;5�_�  �  �          �   o        ����                                                                                                                                                                    
                                                       �                                                                                              o           o           V        ^֣  G �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�   �   �   �            end if;�   �   �   �               end if;�   �   �   �                  end case;�      �   �                     when others =>�   ~   �   �                        end if;�   }      �      (                     bitCounter    := 0;�   |   ~   �      4                     preState      <= waitingSvalid;�   {   }   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   z   |   �      *                     validW(0)     <= '0';�   y   {   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   x   z   �      $               when waitingMready =>�   w   y   �                        end if;�   v   x   �      &                     validW(0) <= '0';�   u   w   �                        else�   t   v   �                           end case;�   s   u   �      &                        when others =>�   r   t   �      !                          end if;�   q   s   �      =                              preState      <= waitingMready;�   p   r   �      3                              s_axis_tready <= '0';�   o   q   �                                  else �   n   p   �      .                              bitCounter := 0;�   m   o   �      0                          if readyW(0) ='1' then�   l   n   �      +                          validW(0) <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      +                          validW(0) <= '0';�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   n   p          1                              bitCounter    := 0;5�_�  �  �          �   n        ����                                                                                                                                                                    
                                                       �                                                                                              n          p          V       ^ٯ     �   m   n          0                          if readyW(0) ='1' then   .                              bitCounter := 0;                               else 5�_�  �  �          �   n        ����                                                                                                                                                                    
                                                       �                                                                                              n          o          V       ^ٱ     �   n   p          =                              preState      <= waitingMready;�   m   o          3                              s_axis_tready <= '0';5�_�  �  �  �      �   m        ����                                                                                                                                                                    
                                                       �                                                                                              m           o           V        ^ٸ     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�      �   �            end if;�   ~   �   �               end if;�   }      �                  end case;�   |   ~   �                     when others =>�   {   }   �                        end if;�   z   |   �      (                     bitCounter    := 0;�   y   {   �      4                     preState      <= waitingSvalid;�   x   z   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   w   y   �      *                     validW(0)     <= '0';�   v   x   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingMready =>�   t   v   �                        end if;�   s   u   �      &                     validW(0) <= '0';�   r   t   �                        else�   q   s   �                           end case;�   p   r   �      &                        when others =>�   o   q   �      !                          end if;�   n   p   �      9                          preState      <= waitingMready;�   m   o   �      /                          s_axis_tready <= '0';�   l   n   �      /                          validW(0)     <= '1';�   k   m   �      !                          end if;�   j   l   �      7                             wirez(0) <= (others=>'0');�   i   k   �                                else �   h   j   �      $                             end if;�   g   i   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   f   h   �      "                             else �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   d   f   �      8                             if s_axis_tdata(7)='1' then�   c   e   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   b   d   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   a   c   �      �                        when 2 =>                                                                           --el y se copia tal cual�   `   b   �      !                          end if;�   _   a   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ^   `   �      -                             inv(0)   <= '0';�   ]   _   �                                else�   \   ^   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   [   ]   �      -                             inv(0)   <= '1';�   Z   \   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   Y   [   �      +                          validW(0) <= '0';�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   l   n          +                          validW(0) <= '1';�   n   p          9                          preState      <= waitingMready;�   m   o          /                          s_axis_tready <= '0';5�_�  �  �          �   t       ����                                                                                                                                                                    
                                                       �                                                                                              m          o          V       ^پ     �   s   t          &                     validW(0) <= '0';5�_�  �  �          �   Z        ����                                                                                                                                                                    
                                                       �                                                                                              Z          Z          V       ^��  H �   Y   Z          +                          validW(0) <= '0';5�_�  �  �          �   o       ����                                                                                                                                                                    
                                                       �                                                                                              Z          Z          V       ^��     �   n   o          !                          end if;5�_�  �  �          �   l        ����                                                                                                                                                                    
                                                       �                                                                                              n          l          V       ^��  I �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �                           end if;�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�      �   �      )   pos_cordic_proc:process (clk) is --{{{�   }      �      %   end process pre_cordic_proc; --}}}�   |   ~   �            end if;�   {   }   �               end if;�   z   |   �                  end case;�   y   {   �                     when others =>�   x   z   �                        end if;�   w   y   �      (                     bitCounter    := 0;�   v   x   �      4                     preState      <= waitingSvalid;�   u   w   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   t   v   �      *                     validW(0)     <= '0';�   s   u   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   r   t   �      $               when waitingMready =>�   q   s   �                        end if;�   p   r   �                        else�   o   q   �                           end case;�   n   p   �      &                        when others =>�   m   o   �      9                          preState      <= waitingMready;�   l   n   �      /                          s_axis_tready <= '0';�   k   m   �      /                          validW(0)     <= '1';�   j   l   �      !                          end if;�   i   k   �      7                             wirez(0) <= (others=>'0');�   h   j   �                                else �   g   i   �      $                             end if;�   f   h   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   e   g   �      "                             else �   d   f   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   c   e   �      8                             if s_axis_tdata(7)='1' then�   b   d   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   a   c   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      �                        when 2 =>                                                                           --el y se copia tal cual�   _   a   �      !                          end if;�   ^   `   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '0';�   \   ^   �                                else�   [   ]   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   Z   \   �      -                             inv(0)   <= '1';�   Y   [   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   X   Z   �      o                        when 1 =>                                                                           --X�   W   Y   �      '                     case bitCounter is�   V   X   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   U   W   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   T   V   �      $               when waitingSvalid =>�   S   U   �                  case preState is�   R   T   �               else�   Q   S   �                  bitCounter    := 0;�   P   R   �      !            inv(0)        <= '0';�   O   Q   �      !            validW(0)     <= '0';�   N   P   �      !            s_axis_tready <= '1';�   M   O   �      +            preState      <= waitingSvalid;�   L   N   �               if rst = '0' then�   K   M   �            if rising_edge(clk) then�   J   L   �         begin�   I   K   �      1      variable bitCounter :integer range 0 to 8 ;�   H   J   �      )   pre_cordic_proc:process (clk) is --{{{�   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   C   E   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   A   C   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   @   B   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   ?   A   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   >   @   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   <   >   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   ;   =   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   :   <   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   9   ;   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   6   8   �      "   signal xyData    : xyDataArray;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   k   m          /                          validW(0)     <= '1';�   m   o          9                          preState      <= waitingMready;�   l   n          /                          s_axis_tready <= '0';5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              n          l          V       ^�k     �   F   H   �       5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              n          l          V       ^�q     �   F   H   �    �   G   H   �    5�_�  �  �          �   G   $    ����                                                                                                                                                                    
                                                       �                                                                                              o          m          V       ^�s     �   F   H   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   G   #    ����                                                                                                                                                                    
                                                       �                                                                                              o          m          V       ^�s     �   F   H   �      $   signal atanLUT : intLUT       :=    X25735.93	15192.80	8027.46	4074.86	2045.34	1023.67	511.96	255.99	128.00	64.00	32.00	16.005�_�  �  �  �      �   G   )    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�{     �   F   H   �      |   signal atanLUT : intLUT       := 25735.93	15192.80	8027.46	4074.86	2045.34	1023.67	511.96	255.99	128.00	64.00	32.00	16.005�_�  �  �          �   G   )    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^ۊ     �   G   I   �         �   G   I   �    5�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^ے     �   G   I   �      7   25736	15193	8027	4075	2045	1024	512	256	128	64	32	165�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^ے     �   G   I   �      7   25736m15193	8027	4075	2045	1024	512	256	128	64	32	165�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^۬     �   G   I   �      7   25736,15193	8027	4075	2045	1024	512	256	128	64	32	165�_�  �  �  �      �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^۴     �   G   I   �      7   25736,15193 8027	4075	2045	1024	512	256	128	64	32	165�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^۶     �   G   I   �      7   25736,15193,8027	4075	2045	1024	512	256	128	64	32	165�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^۸     �   G   I   �      7   25736,15193,8027,4075	2045	1024	512	256	128	64	32	165�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^ۻ     �   G   I   �      7   25736,15193,8027,4075,2045	1024	512	256	128	64	32	165�_�  �             �   H   "    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024	512	256	128	64	32	165�_�  �                H   "    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024.512	256	128	64	32	165�_�                  H   &    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024,512	256	128	64	32	165�_�                 H   *    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024,512,256	128	64	32	165�_�                 H   .    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024,512,256,128	64	32	165�_�                 H   1    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024,512,256,128,64	32	165�_�                 H   4    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   G   I   �      7   25736,15193,8027,4075,2045,1024,512,256,128,64,32	165�_�                 G   $    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      z   signal atanLUT : intLUT       := 25735,	15192.80	8027.46	4074.86	2045.34	1023.67	511.96	255.99	128.00	64.00	32.00	16.005�_�                 G   #    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      $   signal atanLUT : intLUT       :=    7   25736,15193,8027,4075,2045,1024,512,256,128,64,32,165�_�    	             G   $    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      X   signal atanLUT : intLUT       := 25736,15193,8027,4075,2045,1024,512,256,128,64,32,165�_�    
          	   G   Y    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      Y   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64,32,165�_�  	            
   G   S    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      Z   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64,32,16)5�_�  
               G   S    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      Z   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64,32,16)5�_�                 G   T    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      [   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64),32,16)5�_�                 G   T    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��     �   F   H   �      T   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64)5�_�                 F       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^��  J �   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�                 E   Y    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�  K �   D   F   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�                 �        ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�L  M �   �   �   �                              �   �   �   �    5�_�                 �   "    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�l     �   �   �   �      #                        shift_right5�_�               �   "    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�t  N �   �   �   �      "                        shift_righ5�_�                 �   #    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^܁     �   �   �   �      #                        shift_right5�_�                 �        ����                                                                                                                                                                    
                                                       �                                                                                              �           �           V        ^܉     �   �   �   �    �   �   �   �    �   �   �          $                        shift_right(5�_�                 �   2    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ܦ     �   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �    5�_�                 �   =    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ܧ     �   �   �   �      U                        angle <= std_logic_vector(shift_right-signed(wirez(ITER-1)));5�_�                 �   S    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ܭ     �   �   �   �      V                        angle <= std_logic_vector(shift_right(-signed(wirez(ITER-1)));5�_�                 �   S    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ܰ     �   �   �   �      W                        angle <= std_logic_vector(shift_right(-signed(wirez(ITER-1))));5�_�                 G       ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߌ     �   G   J   �         �   G   I   �    5�_�                 H        ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߑ     �   G   I   �    �   H   I   �    5�_�                 H   %    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߓ     �   G   I   �      U   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�                 H   $    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߔ     �   G   I   �      %   signal atanLUT : intLUT       := (    5�_�                 H   %    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߔ     �   G   I   �      &   signal atanLUT : intLUT       := (    !   804	475	251	127	64	32	16	8	4	25�_�                  H   )    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߖ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804	475	251	127	64	32	16	8	4	25�_�    !              H   -    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߘ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475	251	127	64	32	16	8	4	25�_�     "          !   H   1    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߙ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251	127	64	32	16	8	4	25�_�  !  #          "   H   5    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߛ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127	64	32	16	8	4	25�_�  "  $          #   H   8    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߜ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64	32	16	8	4	25�_�  #  %          $   H   ;    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߝ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64,32	16	8	4	25�_�  $  &          %   H   >    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߞ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16	8	4	25�_�  %  '          &   H   @    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߞ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8	4	25�_�  &  (          '   H   B    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߟ     �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4	25�_�  '  )          (   H   D    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߠ  O �   G   I   �      D   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,25�_�  (  *          )   G        ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^ߤ  P �   F   H   �      U   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�  )  +          *   �   X    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^߶  S �   �   �   �      Z                        angle <= std_logic_vector(shift_right(-signed(wirez(ITER-1),8))));5�_�  *  ,          +   �   ,    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^��     �   �   �   �    5�_�  +  -          ,   �       ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^��  T �   �   �   �            �   �   �   �    5�_�  ,  .          -   �       ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^��     �   �   �   �            variable test : signed ;5�_�  -  /          .   �   /    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^�     �   �   �   �      4      variable test : signed range -2**N to 2**N-1);5�_�  .  0          /   �   '    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^�     �   �   �   �      5      variable test : signed range -2**N to 2**(N-1);5�_�  /  1          0   �   )    ����                                                                                                                                                                    
                                                       �                                                                                              �   =       �   G       v   G    ^�
  U �   �   �   �      6      variable test : signed range -2**(N to 2**(N-1);5�_�  0  2          1   �        ����                                                                                                                                                                    
                                                       �                                                                                              �           �           V        ^�2     �   �   �   �    �   �   �   �    �   �   �          9      variable test : signed range -2**(N-1) to 2**(N-1);5�_�  1  3          2   �       ����                                                                                                                                                                    
                                                       �                                                                                              �           �   /       V        ^�3  V �   �   �   �      0      variable y_signed : signed (N-1 downto 0);5�_�  2  4          3   �        ����                                                                                                                                                                    
                                                       �                                                                                              �           �   /       V        ^�9     �   �   �   �       5�_�  3  5          4   �   5    ����                                                                                                                                                                    
                                                       �                                                                                              �           �   /       V        ^�K  W �   �   �   �      6                        test := -signed(wirez(ITER-1);5�_�  4  6          5   �   2    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�U     �   �   �   �      Y                        angle <= std_logic_vector(shift_right(-signed(wirez(ITER-1),8)));5�_�  5  7          6   �   G    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�V     �   �   �   �      M                        angle <= std_logic_vector(-signed(wirez(ITER-1),8)));5�_�  6  8          7   �   G    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�V     �   �   �   �      L                        angle <= std_logic_vector(-signed(wirez(ITER-1)8)));5�_�  7  9          8   �   G    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�W  X �   �   �   �      K                        angle <= std_logic_vector(-signed(wirez(ITER-1))));5�_�  8  :          9   �       ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�h  Y �   �   �          Z                        m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));5�_�  9  ;          :   �       ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�m     �   �   �   �                              �   �   �   �    5�_�  :  <          ;   �   *    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^��  Z �   �   �   �      *                        test := shit_left(5�_�  ;  =          <   �   %    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�  [ �   �   �   �      2                        test := shit_left(test,2);5�_�  <  >          =   �   #    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�     �   �   �   �      3                        test := shit_right(test,2);5�_�  =  ?          >   �   &    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�     �   �   �   �      4                        test := shift_right(test,2);5�_�  >  @          ?   �   &    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�  \ �   �   �   �      3                        test := shift_left(test,2);5�_�  ?  A          @   �   ,    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^�     �   �   �   �                              �   �   �   �    5�_�  @  B          A   �       ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^��  ] �   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));5�_�  A  D          B   �   !    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^��     �   �   �   �      &                        angle <= test;5�_�  B  E  C      D   �   6    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^��  ^ �   �   �   �      7                        angle <= std_logic_vector(test;5�_�  D  F          E   �        ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^��     �   �   �   �    �   �   �   �    5�_�  E  G          F   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^��  _ �   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  F  H          G   �   1    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�     �   �   �   �      4                        test := shift_right(test,2);5�_�  G  I          H   �   1    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�     �   �   �   �      4                        test := shift_right(test,2);5�_�  H  J          I   �   1    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�  ` �   �   �   �      5                        test := shift_right(test,10);5�_�  I  K          J   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�9     �   �   �   �      5                        test := shift_right(test,10);5�_�  J  L          K   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�@  a �   �   �   �      5                        test := shift_right(test,10);5�_�  K  M          L   F       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�j     �   E   G   �      X   --signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  L  N          M   F       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�k     �   E   G   �      W   -signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  M  O          N   H       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�n  b �   G   I   �      F   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  N  P          O   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�;     �   �   �   �      ,      variable test : signed (N-1 downto 0);5�_�  O  Q          P   �   %    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�A     �   �   �   �      3      variable test : signed (-60000 N-1 downto 0);5�_�  P  R          Q   �   %    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�A     �   �   �   �      2      variable test : signed (-60000 -1 downto 0);5�_�  Q  S          R   �   %    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�A     �   �   �   �      1      variable test : signed (-60000 1 downto 0);5�_�  R  T          S   �   %    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�A     �   �   �   �      0      variable test : signed (-60000  downto 0);5�_�  S  U          T   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�D     �   �   �   �      /      variable test : signed (-60000 downto 0);5�_�  T  X          U   �   ,    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�H  c �   �   �   �      /      variable test : signed (-32768 downto 0);5�_�  U  Y  V      X   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�     �   �   �   �      7                        test := -signed(wirez(ITER-1));5�_�  X  Z          Y   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�  e �   �   �   �      7                        test := -signed(wirez(ITER-1));5�_�  Y  [          Z   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^��     �   �   �   �      8                        angle <= std_logic_vector(test);5�_�  Z  \          [   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^��  f �   �   �   �      8                        angle <= std_logic_vector(test);5�_�  [  ]          \   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �                 ^��     �   �   �   �      9                        --test := -signed(wirez(ITER-1));   7                        --test := shift_right(test,10);5�_�  \  ^          ]   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �                 ^��  g �   �   �   �      9                        --test := -signed(wirez(ITER-1));   7                        --test := shift_right(test,10);5�_�  ]  _          ^   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �                 ^��     �   �   �   �      5                        test := shift_right(test,10);�   �   �   �      7                        test := -signed(wirez(ITER-1));5�_�  ^  `          _   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �                 ^��     �   �   �   �      5                        test := shift_right(test,10);5�_�  _  a          `   �        ����                                                                                                                                                                    
                                                       �                                                                                              �          �                 ^��  h �   �   �   �      7                        test := -signed(wirez(ITER-1));5�_�  `  b          a   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��  i �   �   �   �      3      variable test : signed (-32768 downto 32767);5�_�  a  c          b   �        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   �   �   �      6                        test := signed(wirez(ITER-1));5�_�  b  d          c   �   +    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�      �   �   �   �      :                        test := to_integer(wirez(ITER-1));5�_�  c  e          d   �   ?    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�#  j �   �   �   �      A                        test := to_integer(signed(wirez(ITER-1));5�_�  d  f          e   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�.     �   �   �   �      7                        --test := shift_right(test,10);5�_�  e  g          f   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�.  k �   �   �   �      6                        -test := shift_right(test,10);5�_�  f  h          g   �   +    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�?     �   �   �   �      B                        test := to_integer(signed(wirez(ITER-1)));5�_�  g  i          h   �   K    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�F     �   �   �   �      N                        test := to_integer(shift_right(signed(wirez(ITER-1)));5�_�  h  j          i   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�J  l �   �   �   �      5                        test := shift_right(test,10);5�_�  i  k          j   �   L    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�S  m �   �   �   �      O                        test := to_integer(shift_right(signed(wirez(ITER-1))));5�_�  j  l          k   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�\     �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),2));5�_�  k  m          l   �   O    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�]     �   �   �   �      S                        test := to_integer(shift_right(signed(wirez(ITER-1)),102));5�_�  l  n          m   �   8    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�a     �   �   �   �    �   �   �   �    5�_�  m  o          n   �   7    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�d  n �   �   �   �      R                        test := to_integer(shift_right(signed(wirez(ITER-1)),10));5�_�  n  p          o   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�l     �   �   �   �      :                        --angle <= std_logic_vector(test);5�_�  o  q          p   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�l  o �   �   �   �      9                        -angle <= std_logic_vector(test);5�_�  p  r          q   �   2    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�{     �   �   �   �      8                        angle <= std_logic_vector(test);5�_�  q  s          r   �   @    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  p �   �   �   �      B                        angle <= std_logic_vector(to_signed(test);5�_�  r  t          s   �   @    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  q �   �   �   �      C                        angle <= std_logic_vector(to_signed(test));5�_�  s  u          t   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  r �   �   �   �    �   �   �   �    5�_�  t  v          u   f   G    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   e   g   �    �   f   g   �    5�_�  u  w          v   f        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  v  x          w   g   G    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   f   h   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  w  y          x   i   H    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j   �    �   i   j   �    5�_�  x  z          y   i        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  y  �          z   j   H    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��  u �   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  z  �  {      �   F       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   G   I   �      H  -- signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��  v �   G   I   �      G  - signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   �   N    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   �   �   �      S                        test := to_integer(shift_right(-signed(wirez(ITER-1)),10));5�_�  �  �          �   �   O    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   �   �   �      T                        test := to_integer(shift_right(-signed(wirez(ITER-1)),810));5�_�  �  �          �   �   O    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   �   �   �      S                        test := to_integer(shift_right(-signed(wirez(ITER-1)),80));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  w �   �   �   �      R                        test := to_integer(shift_right(signed(wirez(ITER-1)),10));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  x �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),0));5�_�  �  �          �   �   N    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�D     �   �   �   �      R                        test := to_integer(shift_right(-signed(wirez(ITER-1)),8));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�F  y �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),8));5�_�  �  �          �   �   N    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�X     �   �   �   �      R                        test := to_integer(shift_right(-signed(wirez(ITER-1)),1));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�Z  z �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),1));5�_�  �  �          �   �   N    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�l     �   �   �   �      R                        test := to_integer(shift_right(-signed(wirez(ITER-1)),2));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�o  { �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),2));5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   F   H   �      W--   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   F   H   �      V-   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�  �  �          �   H        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  | �   G   I   �      F   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   F   H   �      U   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�  �  �          �   F       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   E   G   �      X   --signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   F       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   E   G   �      W   -signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   i       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j   �      b                                --wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   i       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j   �      a                               --wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   i       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j   �      `                               -wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   i       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   h   j          _                               wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   j        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   j   l   �    5�_�  �  �          �   j        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   i   k   �      _                                wirez(0) <= std_logic_vector(to_signed(-3217,wirez(0)'length));5�_�  �  �          �   k        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   j   k           5�_�  �  �          �   f        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   e   g   �      a                                --wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  �  �          �   f        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   e   g   �      `                                -wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  �  �          �   g        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��  } �   f   h   �      ^                                wirez(0) <= std_logic_vector(to_signed(3217,wirez(0)'length));5�_�  �  �  �      �   H        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   G   I   �      H--   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   H        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   G   I   �      G-   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   F        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  ~ �   E   G   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   H       ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�)   �   H   J   �         �   H   J   �    5�_�  �  �          �   I        ����                                                                                                                                                                    
                                                       �                                                                                              I          I          V       ^�>     �   H   I             constant SCALE := 1024;5�_�  �  �          �   2        ����                                                                                                                                                                    
                                                       �                                                                                              I          I          V       ^�D  � �   1   3   �    �   2   3   �    5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�M  � �   1   3   �         constant SCALE := 1024;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�S  � �   1   3   �      "   constant SCALE := natural 1024;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�Y  � �   1   3   �      $   constant SCALE := natural :=1024;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�`  � �   1   3   �      #   constant SCALE = natural :=1024;5�_�  �  �          �   g   G    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�j     �   f   h   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  �  �          �   j   H    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�m  � �   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�  � �   1   3   �      #   constant SCALE : natural :=1024;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��  � �   1   3   �      "   constant SCALE : natural :=512;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��  � �   1   3   �      "   constant SCALE : natural :=256;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��  � �   1   3   �      "   constant SCALE : natural :=127;5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��     �   1   3   �      !   constant SCALE : natural :=64;5�_�  �  �          �   2   !    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��     �   1   3   �      #   constant SCALE : natural :=1025;5�_�  �  �          �   �   N    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��     �   �   �   �      R                        test := to_integer(shift_right(-signed(wirez(ITER-1)),4));5�_�  �  �          �   �   M    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��  � �   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),4));5�_�  �  �  �      �   J       ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^��     �   I   K   �         �   I   K   �    5�_�  �  �          �   I   '    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   H   J   �    �   I   J   �    5�_�  �  �          �   J   %    ����                                                                                                                                                                    
                                                       �                                                                                              L          L          V       ^��     �   I   K   �      F   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   J   $    ����                                                                                                                                                                    
                                                       �                                                                                              L          L          V       ^��     �   I   K   �      %   signal atanLUT : intLUT       := (       512	302	160	81	41	20	10	5	3	15�_�  �  �          �   J   )    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512	302	160	81	41	20	10	5	3	15�_�  �  �          �   J   -    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302	160	81	41	20	10	5	3	15�_�  �  �          �   J   1    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160	81	41	20	10	5	3	15�_�  �  �          �   J   4    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81	41	20	10	5	3	15�_�  �  �          �   J   7    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41	20	10	5	3	15�_�  �  �          �   J   :    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41,20	10	5	3	15�_�  �  �          �   J   =    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10	5	3	15�_�  �  �          �   J   ?    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5	3	15�_�  �  �          �   J   A    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3	15�_�  �  �          �   J   C    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      C   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,15�_�  �  �          �   J   D    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      E   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);5�_�  �  �          �   J   D    ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   I   K   �      E   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1)l5�_�  �  �          �   I        ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��     �   H   J   �      F   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              K          K          V       ^��  � �   1   3   �      #   constant SCALE : natural :=1023;5�_�  �  �  �      �   F   \    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^��     �   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**N  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   F   ^    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^��  � �   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**16N  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..5�_�  �  �          �   �   6    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);5�_�  �  �          �   �   6    ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^�.     �   �   �   �      B                        m_axis_tdata <= wirez(ITER-1)(N downto 7);5�_�  �  �          �   �   ?    ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^�0  � �   �   �   �      B                        m_axis_tdata <= wirez(ITER-1)(7 downto 7);5�_�  �  �          �   �   O    ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^�B     �   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));5�_�  �  �          �   �   X    ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^�D  � �   �   �   �      ]                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(7 downto 7)));5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^��     �   F   H   �      X--   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^��     �   F   H   �      W-   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);5�_�  �  �          �   J        ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^��     �   I   K   �      E   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);5�_�  �  �          �   2       ����                                                                                                                                                                    
                                                       �                                                                                              �   5       �   ;       v   ;    ^��  � �   1   3   �      #   constant SCALE : natural :=2047;5�_�  �  �  �      �   i        ����                                                                                                                                                                                                                            �                                                                                              f          o                 ^�     �   h   i          `                                --wirez(0) <= std_logic_vector(to_signed(3217,wirez(0)'length));5�_�  �  �          �   k       ����                                                                                                                                                                                                                            �                                                                                              f          n                 ^�  � �   j   k          a                                --wirez(0) <= std_logic_vector(to_signed(-3217,wirez(0)'length));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   3       �   3       V   3    ^��     �   �   �   �      L                        --angle <= std_logic_vector(-signed(wirez(ITER-1)));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   3       �   3       V   3    ^��  � �   �   �   �      K                        -angle <= std_logic_vector(-signed(wirez(ITER-1)));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   3       �   3       V   3    ^��  � �   �   �   �      E                        angle <= std_logic_vector(to_signed(test,N));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   3       �   3       V   3    ^��     �   �   �   �      K                        --angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   3       �   3       V   3    ^��     �   �   �   �      J                        -angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^��  � �   �   �   �      E                        angle <= std_logic_vector(to_signed(test,N));�   �   �   �      Q                        test := to_integer(shift_right(signed(wirez(ITER-1)),0));5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^��     �   �   �   �                              �   �   �   �    5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^      �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^      �   �   �          (                     bitCounter    := 0;5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^ 
     �   �   �   �      +                        bitCounter    := 0;5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^      �   �   �   �      (                        if bitCounter = 5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^ X     �   �   �   �      -                     if(inv(ITER-1)='1') then5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^ Y     �   �   �   �      -                     if inv(ITER-1)='1') then5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^ }     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^      �   �   �   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          v       ^ �     �   �   �   �      G   variable angle     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �          J   variable angleVar     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �          M      variable angleVar     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �            variable test : integer;5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      +      variable test : integer range -2**N ;5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      *      variable test : integer range 2**N ;5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      -      variable test : integer range 2**N)-1 ;5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      .      variable test : integer range *2**N)-1 ;5�_�  �  �          �   �   $    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      .      variable test : integer range )2**N)-1 ;5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      .      variable test : integer range (2**N)-1 ;5�_�  �  �          �   �   *    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      /      variable test : integer range (2**(N)-1 ;5�_�  �  �          �   �   0    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �     �   �   �   �      2      variable test : integer range (2**(N-1))-1 ;5�_�  �  �          �   �   8    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �  � �   �   �   �      B      variable test : integer range (2**(N-1))-1 downto 2**(N-1) ;5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^ �  � �   �   �          0                        if bitCounter = '1' then5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^     �   �   �   �      R                        test := to_integer(shift_right(-signed(wirez(ITER-1)),0));5�_�  �  �          �   �   +    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^     �   �   �   �      G                        test := to_integer((-signed(wirez(ITER-1)),0));5�_�  �             �   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^     �   �   �   �      F                        test := to_integer(-signed(wirez(ITER-1)),0));5�_�  �                �   A    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^     �   �   �   �      E                        test := to_integer(-signed(wirez(ITER-1))0));5�_�                  �   A    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^  � �   �   �   �      D                        test := to_integer(-signed(wirez(ITER-1))));5�_�                 �   2    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^1  � �   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));5�_�                 �   2    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^F     �   �   �   �      T                        angle <= std_logic_vector(test) ; ---signed(wirez(ITER-1)));5�_�                 �   =    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^J  � �   �   �   �      [                        angle <= std_logic_vector(signed(test) ; ---signed(wirez(ITER-1)));5�_�                 �   2    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^P  � �   �   �   �      \                        angle <= std_logic_vector(signed(test)) ; ---signed(wirez(ITER-1)));5�_�                 �   @    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^U  � �   �   �   �      _                        angle <= std_logic_vector(to_signed(test)) ; ---signed(wirez(ITER-1)));5�_�    	           �   A    ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^s     �   �   �   �      b                        angle <= std_logic_vector(to_signed(test,16)) ; ---signed(wirez(ITER-1)));5�_�    
          	   �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�  � �   �   �   �      a                        angle <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�  	            
   �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�     �   �   �   �    �   �   �   �    5�_�  
               �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�     �   �   �   �                              �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�     �   �   �   �                              �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�     �   �   �                               else5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   A       �   B       v   B    ^�     �   �   �   �      ]                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(7 downto 0)));5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^�     �   �   �   �      B                        m_axis_tdata <= wirez(ITER-1)(7 downto 0);�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^�  � �   �   �                               end if;5�_�                 �   +    ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^�  � �   �   �   �      C                        test := to_integer(-signed(wirez(ITER-1)));5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^     �   �   �   �      D                        --m_axis_tdata <= wirez(ITER-1)(7 downto 0);5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �          �                 ^     �   �   �   �      C                        -m_axis_tdata <= wirez(ITER-1)(7 downto 0);5�_�                 �   (    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^
     �   �   �   �      B                        m_axis_tdata <= wirez(ITER-1)(7 downto 0);�   �   �   �    5�_�                 �   K    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^     �   �   �   �      e                        m_axis_tdata <= std_logic_vector(to_signed(test,N))wirez(ITER-1)(7 downto 0);5�_�                 �   (    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^     �   �   �   �      K                        m_axis_tdata <= std_logic_vector(to_signed(test,N))5�_�                 �   (    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^     �   �   �   �      (                        m_axis_tdata <= 5�_�                 �   (    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^*  � �   �   �   �      B                                        wirez(ITER-1)(7 downto 0);5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^D     �   �   �   �    �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^E     �   �   �   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^J     �   �   �   �      H      signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^N  � �   �   �   �      J      variable angle     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^Z     �   �   �   �    �   �   �   �    5�_�                 �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^\     �   �   �   �      h                        angle        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�                  �   &    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^^     �   �   �   �      k                        angleVar        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�    !              �   %    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^_     �   �   �   �      j                        angleVar       <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�     "          !   �   %    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^_     �   �   �   �      i                        angleVar      <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�  !  #          "   �   %    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^c     �   �   �   �    �   �   �   �    5�_�  "  %          #   �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^d     �   �   �   �      C                        test := to_integer(-signed(wirez(ITER-1)));5�_�  #  &  $      %   �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^o     �   �   �   �      C                        anle := to_integer(-signed(wirez(ITER-1)));5�_�  %  )          &   �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^q     �   �   �   �      D                        angle := to_integer(-signed(wirez(ITER-1)));5�_�  &  *  (      )   �   $    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^�     �   �   �   �      G                        angleVar := to_integer(-signed(wirez(ITER-1)));�   �   �   �    5�_�  )  +          *   �   G    ����                                                                                                                                                                                                                            �                                                                                              �   G       �   h       v   h    ^�     �   �   �   �      j                        angleVar := std_logic_vector(to_signed(test,N))to_integer(-signed(wirez(ITER-1)));5�_�  *  ,          +   �   ?    ����                                                                                                                                                                                                                            �                                                                                              �   ?       �   B       v   B    ^�  � �   �   �   �      H                        angleVar := std_logic_vector(to_signed(test,N));�   �   �   �    5�_�  +  -          ,   �       ����                                                                                                                                                                                                                            �                                                                                              �   ?       �   `       v   B    ^�  � �   �   �          h                        angleVar     <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�  ,  /          -   �       ����                                                                                                                                                                                                                            �                                                                                              �   ?       �   `       v   B    ^�  � �   �   �          9                        m_axis_tdata <= test(7 downto 0);5�_�  -  0  .      /   �        ����                                                                                                                                                                                                                            �                                                                                              �   *       �   *       V   *    ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      +                        bitCounter    := 0;�   �   �   �      8                        bitCounter    := bitCounter + 1;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �      D                                        --wirez(ITER-1)(7 downto 0);�   �   �   �      K                        --angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �      :                       -- angle <= std_logic_vector(test);�   �   �   �      7                        --test := shift_right(test,10);�   �   �   �      G                        --angle <= std_logic_vector(to_signed(test,N));�   �   �   �      S                        --test := to_integer(shift_right(signed(wirez(ITER-1)),0));�   �   �   �      _                        --m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(7 downto 0)));�   �   �   �      h                        angle        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));�   �   �   �      G                        --angle <= std_logic_vector(to_signed(test,N));�   �   �   �      7                        --test := shift_right(test,10);�   �   �   �      9                        --test := -signed(wirez(ITER-1));�   �   �   �                           end if;�   �   �   �      B                        test := to_integer(signed(wirez(ITER-1)));�   �   �   �                           else�   �   �   �      f                        angleVar := std_logic_vector(to_signed(to_integer(-signed(wirez(ITER-1))),N));�   �   �   �      G                        test     := to_integer(-signed(wirez(ITER-1)));�   �   �   �      -                     if inv(ITER-1)='1'  then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      M      variable angleVar     : std_logic_vector(N-1 downto 0):= (others=>'0');�   �   �   �      C      variable test : integer range (2**(N-1))-1 downto -2**(N-1) ;�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�      �   �            end if;�   ~   �   �               end if;�   }      �                  end case;�   |   ~   �                     when others =>�   {   }   �                        end if;�   z   |   �      (                     bitCounter    := 0;�   y   {   �      4                     preState      <= waitingSvalid;�   x   z   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   w   y   �      *                     validW(0)     <= '0';�   v   x   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingMready =>�   t   v   �                        end if;�   s   u   �                        else�   r   t   �                           end case;�   q   s   �      &                        when others =>�   p   r   �      9                          preState      <= waitingMready;�   o   q   �      /                          s_axis_tready <= '0';�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      7                             wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   d   f   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   c   e   �      �                        when 2 =>                                                                           --el y se copia tal cual�   b   d   �      !                          end if;�   a   c   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   [   ]   �      o                        when 1 =>                                                                           --X�   Z   \   �      '                     case bitCounter is�   Y   [   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   X   Z   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case preState is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      !            inv(0)        <= '0';�   R   T   �      !            validW(0)     <= '0';�   Q   S   �      !            s_axis_tready <= '1';�   P   R   �      +            preState      <= waitingSvalid;�   O   Q   �               if rst = '0' then�   N   P   �            if rising_edge(clk) then�   M   O   �         begin�   L   N   �      1      variable bitCounter :integer range 0 to 8 ;�   K   M   �      )   pre_cordic_proc:process (clk) is --{{{�   I   K   �      G--   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);�   H   J   �      H--   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);�   G   I   �      W--   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);�   F   H   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**16  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   D   F   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   B   D   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   A   C   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   @   B   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   ?   A   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   ;   =   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   :   <   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   8   :   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal posState  : axiStates := waitingSvalid;�   4   6   �      1   signal preState  : axiStates := waitingSvalid;�   3   5   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   2   4   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �      $   constant SCALE : natural :=18000;�   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          C                        test := to_integer(-signed(wirez(ITER-1)));�   �   �          f                        angleVar := std_logic_vector(to_signed(to_integer(-signed(wirez(ITER-1))),N));5�_�  /  1          0   �   9    ����                                                                                                                                                                                                                            �                                                                                              �   *       �   *       V   *    ^2     �   �   �   �    �   �   �   �    5�_�  0  2          1   �       ����                                                                                                                                                                                                                            �                                                                                              �   *       �   *       V   *    ^3     �   �   �   �      h                        angle        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�  1  3          2   �   9    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^A     �   �   �   �      h                        angle        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));�   �   �   �    5�_�  2  4          3   �   F    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^C     �   �   �   �      u                        angle        <= std_logic_vector(wirez(ITER-1)to_signed(test,N)) ; ---signed(wirez(ITER-1)));5�_�  3  5          4   �   F    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^C     �   �   �   �      F                        angle        <= std_logic_vector(wirez(ITER-1)5�_�  4  6          5   �   F    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^E     �   �   �   �      G                        angle        <= std_logic_vector(wirez(ITER-1);5�_�  5  7          6   �   9    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^G     �   �   �   �      H                        angle        <= std_logic_vector(wirez(ITER-1));5�_�  6  9          7   �   J    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^L     �   �   �   �      L                        angle        <= std_logic_vector(not)wirez(ITER-1));5�_�  7  :  8      9   �   <    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^~     �   �   �   �      O                        angle        <= std_logic_vector(not)wirez(ITER-1))+1);5�_�  9  ;          :   �   (    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   8       v   8    ^�     �   �   �   �      O                        angle        <= std_logic_vector(not(wirez(ITER-1))+1);5�_�  :  <          ;   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   8       v   8    ^�     �   �   �   �      >                        angle        <= not(wirez(ITER-1))+1);5�_�  ;  =          <   �   M    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   8       v   8    ^�  � �   �   �   �      O                        angle        <= not(wirez(ITER-1))+std_logic_vector(1);5�_�  <  >          =   �   L    ����                                                                                                                                                                                                                            �                                                                                              �   (       �   8       v   8    ^�     �   �   �   �      P                        angle        <= not(wirez(ITER-1))+std_logic_vector(1));5�_�  =  ?          >   �   O    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�     �   �   �   �      S                        angle        <= not(wirez(ITER-1))+std_logic_vector(to_1));5�_�  >  @          ?   �   X    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�  � �   �   �   �      [                        angle        <= not(wirez(ITER-1))+std_logic_vector(to_integer(1));5�_�  ?  A          @   �   Z    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�  � �   �   �   �      \                        angle        <= not(wirez(ITER-1))+std_logic_vector(to_integer(1)));5�_�  @  B          A   �   L    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�     �   �   �   �      [                        angle        <= not(wirez(ITER-1))+std_logic_vector(to_integer(1));5�_�  A  C          B   �   L    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�     �   �   �   �      Z                        angle        <= not(wirez(ITER-1))+std_logic_vector(o_integer(1));5�_�  B  D          C   �   L    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   N       v   N    ^�  � �   �   �   �      Y                        angle        <= not(wirez(ITER-1))+std_logic_vector(_integer(1));5�_�  C  E          D   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �   �      X                        angle        <= not(wirez(ITER-1))+std_logic_vector(integer(1));5�_�  D  F          E   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �   �      @                        angle        <= not(wirez(ITER-1))+l1));5�_�  E  G          F   �   <    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �   �      ?                        angle        <= not(wirez(ITER-1))+1));5�_�  F  H          G   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �   �      >                        angle        <= not(wirez(ITER-1))+1);5�_�  G  I          H   �   =    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�  � �   �   �   �      ?                        angle        <= not(wirez(ITER-1))+"1);5�_�  H  J          I   �   L    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�  � �   �   �   �      N                        angle        <= not(wirez(ITER-1))+"1"&(others=>'0'));5�_�  I  K          J   �       ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �   �    �   �   �   �    5�_�  J  L          K   �       ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^�     �   �   �          G                        test     := to_integer(-signed(wirez(ITER-1)));5�_�  K  M          L   �       ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^#     �   �   �   �      M      variable angleVar     : std_logic_vector(N-1 downto 0):= (others=>'0');5�_�  L  N          M   �   2    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^;     �   �   �   �      C      variable angleVar     : signed(N-1 downto 0):= (others=>'0');5�_�  M  O          N   �   2    ����                                                                                                                                                                                                                            �                                                                                              �   ;       �   S       v   S    ^>  � �   �   �   �      ;      variable angleVar     : signed(N-1 downto 0)rs=>'0');5�_�  N  P          O   �   $    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^I     �   �   �   �      f                        angleVar := std_logic_vector(to_signed(to_integer(-signed(wirez(ITER-1))),N));5�_�  O  Q          P   �   :    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^R  � �   �   �   �      @                        angleVar := -signed(wirez(ITER-1))),N));5�_�  P  R          Q   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^X  � �   �   �          M                        angle        <= not(wirez(ITER-1))+"1"&(others=>'0');5�_�  Q  S          R   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^f  � �   �   �   �    �   �   �   �    5�_�  R  T          S   �   $    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^i  � �   �   �   �      ;                        angleVar := -signed(wirez(ITER-1));5�_�  S  U          T   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^w     �   �   �   �      :                       -- angle <= std_logic_vector(test);5�_�  T  V          U   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^w     �   �   �   �      9                       - angle <= std_logic_vector(test);5�_�  U  W          V   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^w     �   �   �   �      8                        angle <= std_logic_vector(test);5�_�  V  X          W   �   1    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^{  � �   �   �   �      7                       angle <= std_logic_vector(test);5�_�  W  \          X   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �          C      variable test : integer range (2**(N-1))-1 downto -2**(N-1) ;5�_�  X  l  Y      \   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �          B                        test := to_integer(signed(wirez(ITER-1)));5�_�  \  m  ]      l   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �                           �   �   �   �    5�_�  l  n          m   �   9    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�  � �   �   �   �      ;                       angle <= std_logic_vector(angleVar);5�_�  m  o          n   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�  � �   �   �          G                        test     := to_integer(-signed(wirez(ITER-1)));5�_�  n  p          o   �   :    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      B                       angle <= std_logic_vector(angleVar and 12);5�_�  o  q          p   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      D                       angle <= std_logic_vector(angleVar &&and 12);5�_�  p  r          q   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      C                       angle <= std_logic_vector(angleVar &and 12);5�_�  q  s          r   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      B                       angle <= std_logic_vector(angleVar &nd 12);5�_�  r  t          s   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      A                       angle <= std_logic_vector(angleVar &d 12);5�_�  s  u          t   �   :    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      @                       angle <= std_logic_vector(angleVar & 12);5�_�  t  v          u   �   =    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�  � �   �   �   �      C                       angle <= std_logic_vector(angleVar AND& 12);5�_�  u  w          v   �   1    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      B                       angle <= std_logic_vector(angleVar AND 12);5�_�  v  x          w   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      I                       angle <= std_logic_vector("00" & angleVar AND 12);5�_�  w  y          x   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      H                       angle <= std_logic_vector("00" & angleVar ND 12);5�_�  x  z          y   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      G                       angle <= std_logic_vector("00" & angleVar D 12);5�_�  y  {          z   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      F                       angle <= std_logic_vector("00" & angleVar  12);5�_�  z  |          {   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      E                       angle <= std_logic_vector("00" & angleVar 12);5�_�  {  }          |   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      D                       angle <= std_logic_vector("00" & angleVar 2);5�_�  |  ~          }   �   @    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�  � �   �   �   �      C                       angle <= std_logic_vector("00" & angleVar );5�_�  }            ~   �   4    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      B                       angle <= std_logic_vector("00" & angleVar);5�_�  ~  �             �   F    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      H                       angle <= std_logic_vector("00000000" & angleVar);5�_�    �          �   �   P    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      T                       angle <= std_logic_vector("00000000" & angleVar(7 downto 9));5�_�  �  �          �   �   P    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�  � �   �   �   �      T                       angle <= std_logic_vector("00000000" & angleVar(7 downto 9));5�_�  �  �          �   �   1    ����                                                                                                                                                                                                                            �                                                                                              �   1       �   =       v   =    ^�  � �   �   �   �      T                       angle <= std_logic_vector("00000000" & angleVar(7 downto 0));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   1       �   =       v   =    ^
  � �   �   �   �      G                       angle <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   1       �   =       v   =    ^     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   1       �   =       v   =    ^     �   �   �   �      N                       m_axis_tdata <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   1       �   =       v   =    ^#     �   �   �   �      E                       ang <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �   9    ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^)  � �   �   �   �      G                       angle <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^:     �   �   �   �                              �   �   �   �    5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^H     �   �   �   �      (                        if bitCounter = 5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^W     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^X     �   �   �          N                       m_axis_tdata <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �   E    ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^c     �   �   �   �      R                           m_axis_tdata <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �   P    ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^f     �   �   �   �      T                           m_axis_tdata <= std_logic_vector(angleVar(N-1 downto 0));5�_�  �  �          �   �   P    ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^g     �   �   �   �      T                           m_axis_tdata <= std_logic_vector(angleVar(N-1 downto 9));5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �   9       �   D       v   D    ^l     �   �   �   �       5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^s     �   �   �          +                        bitCounter    := 0;   }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato   �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   -                        readyW(ITER)  <= '1';5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^t     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^u     �   �   �          -                        readyW(ITER)  <= '1';�   �   �          �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �          }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �          +                        bitCounter    := 0;5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^{     �   �   �                                  15�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^|     �   �   �           5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �                              �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      *                     m_axis_tvalid <= '1';5�_�  �  �          �   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      *                     m_axis_tvalid <= '-';5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �       5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          s5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          *                     m_axis_tvalid <= '0';5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �                                 �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          .                           bitCounter    := 0;   �                           posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          0                           readyW(ITER)  <= '1';5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �           5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �    5�_�  �  �          �   �   -    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  �  �          �   �   -    ����                                                                                                                                                                                                                            �                                                                                              �   -       �   -       V   -    ^�     �   �   �          K                        --angle <= std_logic_vector(signed(wirez(ITER-1)));   D                                        --wirez(ITER-1)(7 downto 0);5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �       	                              9                        --test := -signed(wirez(ITER-1));   7                        --test := shift_right(test,10);   G                        --angle <= std_logic_vector(to_signed(test,N));   j                        --angle        <= std_logic_vector(to_signed(test,N)) ; ---signed(wirez(ITER-1)));   _                        --m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(7 downto 0)));   S                        --test := to_integer(shift_right(signed(wirez(ITER-1)),0));   G                        --angle <= std_logic_vector(to_signed(test,N));   7                        --test := shift_right(test,10);5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �          ;                       angle <= std_logic_vector(angleVar);�   �   �          N                       m_axis_tdata <= std_logic_vector(angleVar(7 downto 0));5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        m_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �                              end if�   �   �   �      0                           readyW(ITER)  <= '1';�   �   �   �      �                           posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �                              else�   �   �   �      T                           m_axis_tdata <= std_logic_vector(angleVar(N-1 downto 8));�   �   �   �      �                           m_axis_tvalid <= '1';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      0                        if bitCounter = '1' then�   �   �   �      8                        bitCounter    := bitCounter + 1;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �      A                     angle         <= std_logic_vector(angleVar);�   �   �   �      M                     m_axis_tdata  <= std_logic_vector(angleVar(7 downto 0));�   �   �   �                           end if;�   �   �   �      :                        angleVar := signed(wirez(ITER-1));�   �   �   �                           else�   �   �   �      ;                        angleVar := -signed(wirez(ITER-1));�   �   �   �      -                     if inv(ITER-1)='1'  then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      3      variable angleVar     : signed(N-1 downto 0);�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�      �   �            end if;�   ~   �   �               end if;�   }      �                  end case;�   |   ~   �                     when others =>�   {   }   �                        end if;�   z   |   �      (                     bitCounter    := 0;�   y   {   �      4                     preState      <= waitingSvalid;�   x   z   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   w   y   �      *                     validW(0)     <= '0';�   v   x   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingMready =>�   t   v   �                        end if;�   s   u   �                        else�   r   t   �                           end case;�   q   s   �      &                        when others =>�   p   r   �      9                          preState      <= waitingMready;�   o   q   �      /                          s_axis_tready <= '0';�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      7                             wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   d   f   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   c   e   �      �                        when 2 =>                                                                           --el y se copia tal cual�   b   d   �      !                          end if;�   a   c   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   [   ]   �      o                        when 1 =>                                                                           --X�   Z   \   �      '                     case bitCounter is�   Y   [   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   X   Z   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case preState is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      !            inv(0)        <= '0';�   R   T   �      !            validW(0)     <= '0';�   Q   S   �      !            s_axis_tready <= '1';�   P   R   �      +            preState      <= waitingSvalid;�   O   Q   �               if rst = '0' then�   N   P   �            if rising_edge(clk) then�   M   O   �         begin�   L   N   �      1      variable bitCounter :integer range 0 to 8 ;�   K   M   �      )   pre_cordic_proc:process (clk) is --{{{�   I   K   �      G--   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);�   H   J   �      H--   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);�   G   I   �      W--   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);�   F   H   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**16  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   D   F   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   B   D   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   A   C   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   @   B   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   ?   A   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   ;   =   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   :   <   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   8   :   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal posState  : axiStates := waitingSvalid;�   4   6   �      1   signal preState  : axiStates := waitingSvalid;�   3   5   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   2   4   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �      $   constant SCALE : natural :=18000;�   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          L                     m_axis_tdata <= std_logic_vector(angleVar(7 downto 0));�   �   �          4                     posState      <= waitingMready;�   �   �          (                     bitCounter    := 0;�   �   �          *                     m_axis_tvalid <= '1';�   �   �          *                     readyW(ITER)  <= '0';�   �   �          9                     angle <= std_logic_vector(angleVar);5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        m_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �                              end if�   �   �   �      0                           readyW(ITER)  <= '1';�   �   �   �      �                           posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �                              else�   �   �   �      U                           m_axis_tdata  <= std_logic_vector(angleVar(N-1 downto 8));�   �   �   �      �                           m_axis_tvalid <= '1';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      0                        if bitCounter = '1' then�   �   �   �      8                        bitCounter    := bitCounter + 1;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �      A                     angle         <= std_logic_vector(angleVar);�   �   �   �      M                     m_axis_tdata  <= std_logic_vector(angleVar(7 downto 0));�   �   �   �                           end if;�   �   �   �      :                        angleVar := signed(wirez(ITER-1));�   �   �   �                           else�   �   �   �      ;                        angleVar := -signed(wirez(ITER-1));�   �   �   �      -                     if inv(ITER-1)='1'  then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      3      variable angleVar     : signed(N-1 downto 0);�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�      �   �            end if;�   ~   �   �               end if;�   }      �                  end case;�   |   ~   �                     when others =>�   {   }   �                        end if;�   z   |   �      (                     bitCounter    := 0;�   y   {   �      4                     preState      <= waitingSvalid;�   x   z   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   w   y   �      *                     validW(0)     <= '0';�   v   x   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingMready =>�   t   v   �                        end if;�   s   u   �                        else�   r   t   �                           end case;�   q   s   �      &                        when others =>�   p   r   �      9                          preState      <= waitingMready;�   o   q   �      /                          s_axis_tready <= '0';�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      7                             wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   d   f   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   c   e   �      �                        when 2 =>                                                                           --el y se copia tal cual�   b   d   �      !                          end if;�   a   c   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   [   ]   �      o                        when 1 =>                                                                           --X�   Z   \   �      '                     case bitCounter is�   Y   [   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   X   Z   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case preState is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      !            inv(0)        <= '0';�   R   T   �      !            validW(0)     <= '0';�   Q   S   �      !            s_axis_tready <= '1';�   P   R   �      +            preState      <= waitingSvalid;�   O   Q   �               if rst = '0' then�   N   P   �            if rising_edge(clk) then�   M   O   �         begin�   L   N   �      1      variable bitCounter :integer range 0 to 8 ;�   K   M   �      )   pre_cordic_proc:process (clk) is --{{{�   I   K   �      G--   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);�   H   J   �      H--   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);�   G   I   �      W--   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);�   F   H   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**16  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   D   F   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   B   D   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   A   C   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   @   B   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   ?   A   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   ;   =   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   :   <   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   8   :   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal posState  : axiStates := waitingSvalid;�   4   6   �      1   signal preState  : axiStates := waitingSvalid;�   3   5   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   2   4   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �      $   constant SCALE : natural :=18000;�   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          �                           m_axis_tvalid <= '1';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �          T                           m_axis_tdata <= std_logic_vector(angleVar(N-1 downto 8));5�_�  �  �          �   �        ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^     �   �   �   �         end generate;�   �   �   �               );�   �   �   �                 rst     => rst�   �   �   �                 clk     => clk,�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �            port  map (�   �   �   �            generic map(N,j)�   �   �   �            iteration: cordic_iter�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �         begin�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �               end if;�   �   �   �                  end if;�   �   �   �                     end case;�   �   �   �                           end if;�   �   �   �      -                        m_axis_tvalid <= '0';�   �   �   �                           else�   �   �   �                              end if�   �   �   �      0                           readyW(ITER)  <= '1';�   �   �   �      �                           posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      .                           bitCounter    := 0;�   �   �   �      �                           m_axis_tvalid <= '0';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �                              else�   �   �   �      U                           m_axis_tdata  <= std_logic_vector(angleVar(N-1 downto 8));�   �   �   �      �                           m_axis_tvalid <= '1';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      0                        if bitCounter = '1' then�   �   �   �      8                        bitCounter    := bitCounter + 1;�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      '                  when waitingMready =>�   �   �   �                        end if;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �      (                     bitCounter    := 0;�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �      A                     angle         <= std_logic_vector(angleVar);�   �   �   �      M                     m_axis_tdata  <= std_logic_vector(angleVar(7 downto 0));�   �   �   �                           end if;�   �   �   �      :                        angleVar := signed(wirez(ITER-1));�   �   �   �                           else�   �   �   �      ;                        angleVar := -signed(wirez(ITER-1));�   �   �   �      -                     if inv(ITER-1)='1'  then�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      $               when waitingSvalid =>�   �   �   �                  case posState is�   �   �   �               else�   �   �   �                  bitCounter := 0;�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �      -            angle         <= (others => '0');�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �               if rst = '0' then�   �   �   �            if rising_edge(clk) then�   �   �   �         begin�   �   �   �      3      variable angleVar     : signed(N-1 downto 0);�   �   �   �      1      variable bitCounter :integer range 0 to 8 ;�   �   �   �      )   pos_cordic_proc:process (clk) is --{{{�   �   �   �      %   end process pre_cordic_proc; --}}}�      �   �            end if;�   ~   �   �               end if;�   }      �                  end case;�   |   ~   �                     when others =>�   {   }   �                        end if;�   z   |   �      (                     bitCounter    := 0;�   y   {   �      4                     preState      <= waitingSvalid;�   x   z   �      e                     s_axis_tready <= '1';                          --entonces yo tambien estoy listo�   w   y   �      *                     validW(0)     <= '0';�   v   x   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   u   w   �      $               when waitingMready =>�   t   v   �                        end if;�   s   u   �                        else�   r   t   �                           end case;�   q   s   �      &                        when others =>�   p   r   �      9                          preState      <= waitingMready;�   o   q   �      /                          s_axis_tready <= '0';�   n   p   �      /                          validW(0)     <= '1';�   m   o   �      !                          end if;�   l   n   �      7                             wirez(0) <= (others=>'0');�   k   m   �                                else �   j   l   �      $                             end if;�   i   k   �      `                                wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));�   h   j   �      "                             else �   g   i   �      _                                wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));�   f   h   �      8                             if s_axis_tdata(7)='1' then�   e   g   �      �                          if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   d   f   �      f                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   c   e   �      �                        when 2 =>                                                                           --el y se copia tal cual�   b   d   �      !                          end if;�   a   c   �      i                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),N));�   `   b   �      -                             inv(0)   <= '0';�   _   a   �                                else�   ^   `   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),N));�   ]   _   �      -                             inv(0)   <= '1';�   \   ^   �      �                          if s_axis_tdata(7)='1' then                                                       --corrijo cuadrante si X es negativo y lo informo en inv�   [   ]   �      o                        when 1 =>                                                                           --X�   Z   \   �      '                     case bitCounter is�   Y   [   �      �                     bitCounter := bitCounter + 1;                                                          --espero 2 datos de 8 bits.. primero X luego Y�   X   Z   �      �                  if s_axis_tvalid = '1' then                                                               --espero a que entren datos�   W   Y   �      $               when waitingSvalid =>�   V   X   �                  case preState is�   U   W   �               else�   T   V   �                  bitCounter    := 0;�   S   U   �      !            inv(0)        <= '0';�   R   T   �      !            validW(0)     <= '0';�   Q   S   �      !            s_axis_tready <= '1';�   P   R   �      +            preState      <= waitingSvalid;�   O   Q   �               if rst = '0' then�   N   P   �            if rising_edge(clk) then�   M   O   �         begin�   L   N   �      1      variable bitCounter :integer range 0 to 8 ;�   K   M   �      )   pre_cordic_proc:process (clk) is --{{{�   I   K   �      G--   signal atanLUT : intLUT       := ( 512,302,160,81,41,20,10,5,3,1);�   H   J   �      H--   signal atanLUT : intLUT       := ( 804,475,251,127,64,32,16,8,4,2);�   G   I   �      W--   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);�   F   H   �      V   signal atanLUT : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   E   G   �      �   type   intLUT        is array   ( MAX_ITER-1 downto 0 )of integer          range 0 to 2**16  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   D   F   �      `   --defino una tabla con los angulos tal que su arcotangente da 1/2**N (la magia de don Cordic)�   B   D   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   A   C   �      ]   type   ConnectVector is array   ( ITER downto 0 )      of std_logic_vector (N-1 downto 0);�   @   B   �      8   --tambien desperdicio uno al final, son ITER+1 cables�   ?   A   �      S   --defino los cables de datos para la interconexion de las instancias del cordica�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   ;   =   �      �   -- notar el detalle que tiene ITER+1 cable porque se desperdicia un cable pero permite hacer la logica de intercoinexion en el for-generate sin problemas�   :   <   �      l   --con esta dos lineas defino una sere de cables para interconectar las instancias del pipeline del Cordic�   8   :   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   7   9   �      "   signal xyData    : xyDataArray;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   5   7   �      1   signal posState  : axiStates := waitingSvalid;�   4   6   �      1   signal preState  : axiStates := waitingSvalid;�   3   5   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   2   4   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   1   3   �      $   constant SCALE : natural :=18000;�   /   1   �         end component; --}}}�   .   0   �      )          rst           : in  STD_LOGIC);�   -   /   �      (          clk           : in  STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   )   +   �      "          s_valid : in  STD_LOGIC;�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   #   %   �      "          m_ready : in  STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   !   #   �      "          m_valid : out STD_LOGIC;�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�         �            port(�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �      9             N     : natural := 16; --Ancho de la palabra�         �            generic(�         �      !   component cordic_iter is --{{{�         �      )          rst           : in  STD_LOGIC);�         �      (          clk           : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          m_axis_tready : in  STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�   
      �      (          m_axis_tvalid : out STD_LOGIC;�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�      
   �         Port(�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�         �      9             N     : natural := 16; --Ancho de la palabra�         �         generic(�   �   �          �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �          �                           posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �          .                           bitCounter    := 0;�   �   �          0                           readyW(ITER)  <= '1';5�_�  �  �          �   �   0    ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^  � �   �   �   �      �                           m_axis_tvalid <= '0';--y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar5�_�  �  �          �   �       ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^  � �   �   �   �                              end if5�_�  �  �          �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^'     �   �   �   �      0                        if bitCounter = '1' then5�_�  �  �          �   �   )    ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^(     �   �   �   �      /                        if bitCounter = 1' then5�_�  �              �   �   (    ����                                                                                                                                                                                                                            �                                                                                              �           �           V        ^)  � �   �   �   �      .                        if bitCounter = 1 then5�_�  \  ^      l  ]   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �        5�_�  ]  _          ^   �        ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �        5�_�  ^  `          _   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      J                       --angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  _  a          `   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      I                       -angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  `  b          a   �       ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      Y                       m_axis_tdata <= -angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  a  c          b   �   (    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      X                       m_axis_tdata <= -ngle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  b  d          c   �   (    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      Y                       m_axis_tdata <= -angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  c  e          d   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      X                       m_axis_tdata <= angle <= std_logic_vector(signed(wirez(ITER-1)));5�_�  d  f          e   �   ,    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      j                       m_axis_tdata <= angleVar(N-1 downto 8); <= std_logic_vector(signed(wirez(ITER-1)));5�_�  e  g          f   �   >    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�  � �   �   �   �      >                       m_axis_tdata <= angleVar(N-1 downto 8);5�_�  f  h          g   �   '    ����                                                                                                                                                                                                                            �                                                                                              �          �          V       ^�     �   �   �   �      O                       m_axis_tdata <= std_logic_vector(angleVar(N-1 downto 8);5�_�  g  i          h   �   @    ����                                                                                                                                                                                                                            �                                                                                              �   A       �   N       v   N    ^�  � �   �   �   �      P                       m_axis_tdata <= std_logic_vector(angleVar)(N-1 downto 8);5�_�  h  j          i   �   A    ����                                                                                                                                                                                                                            �                                                                                              �   A       �   N       v   N    ^�  � �   �   �   �      B                       m_axis_tdata <= std_logic_vector(angleVar);5�_�  i  k          j   �   @    ����                                                                                                                                                                                                                            �                                                                                              �   A       �   N       v   N    ^"     �   �   �   �      C                       m_axis_tdata <= std_logic_vector(angleVar));5�_�  j              k   �   ;    ����                                                                                                                                                                                                                            �                                                                                              �   A       �   N       v   N    ^#     �   �   �   �      <                       angle <= std_logic_vector(angleVar);(5�_�  X  Z      \  Y   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      2      variable anglear     : signed(N-1 downto 0);5�_�  Y  [          Z   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      1      variable angler     : signed(N-1 downto 0);5�_�  Z              [   �       ����                                                                                                                                                                                                                            �                                                                                              �   $       �   I       v   I    ^�     �   �   �   �      0      variable angle     : signed(N-1 downto 0);5�_�  7          9  8   �   H    ����                                                                                                                                                                                                                            �                                                                                              �   @       �   L       v   L    ^[     �   �   �   �       5�_�  -          /  .   �   *    ����                                                                                                                                                                                                                            �                                                                                              �   *       �   *       V   *    ^�     �   �   �   �      Ceeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   feeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  &      '  )  (   �        ����                                                                                                                                                                                                                            �                                                                                              �           �   "       V   $    ^�     �   �   �        �   �   �   �    �   �   �   �      #std_logic_vector(to_signed(test,N))5�_�  &          (  '   �   $    ����                                                                                                                                                                                                                            �                                                                                              �   $       �   7       v   7    ^�     �   �   �   �      3                        angleVar := irez(ITER-1)));5�_�  #          %  $   �       ����                                                                                                                                                                                                                            �                                                                                              �   (       �   J       v   J    ^j     �   �   �   �      E                        testjh := to_integer(-signed(wirez(ITER-1)));5�_�                 �   B    ����                                                                                                                                                                                                                            �                                                                                              �   +       �   5       v   5    ^c  � �   �   �   �      b                        angle <= std_logic_vector(to_signed(test,10)) ; ---signed(wirez(ITER-1)));5�_�  �  �      �  �   f       ����                                                                                                                                                                                                                            �                                                                                                                               ^��     �   f   g   �    �   e   f   �      7                             wirez(0) <= (others=>'0');5�_�  �  �          �   g       ����                                                                                                                                                                                                                            �                                                                                              g          p                 ^��     �   f   h   �      �                          00if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z�   g   q   �   	   :                          00   if s_axis_tdata(7)='1' then   a                          00      wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));   b                          00      --wirez(0) <= std_logic_vector(to_signed(3217,wirez(0)'length));   $                          00   else    b                          00      wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));   c                          00      --wirez(0) <= std_logic_vector(to_signed(-3217,wirez(0)'length));   &                          00   end if;   !                          00else    9                          00   wirez(0) <= (others=>'0');5�_�  �  �          �   g       ����                                                                                                                                                                                                                            �                                                                                              g          p                 ^��     �   f   q   �   
   �                          --if inv(0)='1' then                                                                --si hay cambio de cuadrante aprovecho para sumarle un offset del angulo al Z   :                          --   if s_axis_tdata(7)='1' then   a                          --      wirez(0) <= std_logic_vector(to_signed(SCALE,wirez(0)'length));   b                          --      --wirez(0) <= std_logic_vector(to_signed(3217,wirez(0)'length));   $                          --   else    b                          --      wirez(0) <= std_logic_vector(to_signed(-SCALE,wirez(0)'length));   c                          --      --wirez(0) <= std_logic_vector(to_signed(-3217,wirez(0)'length));   &                          --   end if;   !                          --else    9                          --   wirez(0) <= (others=>'0');5�_�  �  �          �   f       ����                                                                                                                                                                                                                            �                                                                                              g          p                 ^��     �   e   g          4                          wirez(0) <= (others=>'0');5�_�  �              �   q       ����                                                                                                                                                                                                                            �                                                                                              g          p                 ^��     �   p   r   �      #                          --end if;5�_�  �  �      �  �   _   :    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   ^   `   �      V                             wirex(0) <= std_logic_vector((-signed(s_axis_tdata)),N));5�_�  �  �  �      �   _   Q    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   ^   `   �      U                             wirex(0) <= std_logic_vector((-signed(s_axis_tdata))N));5�_�  �  �          �   _   Q    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   ^   `   �      T                             wirex(0) <= std_logic_vector((-signed(s_axis_tdata))));5�_�  �              �   _   R    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�  � �   ^   `   �      S                             wirex(0) <= std_logic_vector((-signed(s_axis_tdata)));5�_�  �  �      �  �   _   R    ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   ^   `   �      U                             wirex(0) <= std_logic_vector((-signed(s_axis_tdata)),));5�_�  �              �   _       ����                                                                                                                                                                    
                                                       �                                                                                              _   :       _   M       v   M    ^�     �   ^   `        5�_�  �  �      �  �   �   7    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�      �   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(12 downto 7);5�_�  �              �   �   @    ����                                                                                                                                                                    
                                                       �                                                                                              J          J          V       ^�&     �   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(12 downto 5);5�_�  �          �  �   G        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^��     �   F   H   �      V-   signal atanLUT : intLUT       := (25736,15193,8027,4075,2045,1024,512,256,128,64);5�_�  z  |      �  {   i        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   h   j   �      a                                -wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  {  }          |   i        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   h   j   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));5�_�  |  ~          }   j        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   i   k   �      a                                --wirez(0) <= std_logic_vector(to_signed(-3217,wirez(0)'length));5�_�  }            ~   f        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   e   g   �      `                                -wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�  ~  �             f        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�     �   e   g   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));5�_�                �   g        ����                                                                                                                                                                    
                                                       �                                                                                              �          �   1       v   1    ^�  t �   f   h   �      `                                --wirez(0) <= std_logic_vector(to_signed(3217,wirez(0)'length));5�_�  U  W      X  V   �       ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�k     �   �   �   �      3      variable test : signed (-60000 downto 32767);5�_�  V              W   �   ,    ����                                                                                                                                                                    
                                                       �                                                                                              �          �          V       ^�n  d �   �   �   �      3      variable test : signed (-60000 downto 60000);5�_�  B          D  C   �   5    ����                                                                                                                                                                    
                                                       �                                                                                              �   2       �   =       v   =    ^��     �   �   �   �      8                        angle <= std_logic_vector(tes)t;5�_�                 �   "    ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^�m     �   �   �   �      #                        shift_right    5�_�  �          �  �   H       ����                                                                                                                                                                    
                                                       �                                                                                              G   )       G   +       v   +    ^ۯ     �   G   I   �      7   25736,151 3 8027	4075	2045	1024	512	256	128	64	32	165�_�  �          �  �   G   $    ����                                                                                                                                                                    
                                                       �                                                                                              n          l          V       ^�v     �   F   H   �      |   signal atanLUT : intLUT       := e5735.93	15192.80	8027.46	4074.86	2045.34	1023.67	511.96	255.99	128.00	64.00	32.00	16.005�_�  �          �  �   m        ����                                                                                                                                                                    
                                                       �                                                                                              m          o          V       ^ٳ     �   l   p   �      +eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   /eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   9eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �          �  �   q        ����                                                                                                                                                                    
                                                       �                                                                                              q          r          V       ^ր     �   p   s   �      3eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   8eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �  �      �  �   i        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�9     �   i   j   �    �   h   i   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   i       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�:     �   h   j          v                          if readyW(0) = '1' then                           --espero e que este listo para enviar algo5�_�  �  �          �   m       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�]     �   m   n   �                           �   m   o   �                        else    5�_�  �  �          �   o        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�_     �   o   p   �    �   o   p   �      /                          validW(0)     <= '1';5�_�  �  �          �   o        ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�`     �   n   p        5�_�  �  �          �   o       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�a     �   n   p          *                     validW(0)     <= '1';5�_�  �  �          �   o   '    ����                                                                                                                                                                >   
                                                       �                                                                                              o   '       o   '       V   '    ^�c     �   n   p   �      *                     validW(0)     <= '0';5�_�  �              �   o        ����                                                                                                                                                                >   
                                                       �                                                                                              o   '       o   '       V   '    ^�e     �   n   p          &                     validW(0) <= '0';�         �         generic(�         �      9             N     : natural := 16; --Ancho de la palabra�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�      
   �         Port(�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   
      �      (          m_axis_tvalid : out STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�         �      (          m_axis_tready : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          clk           : in  STD_LOGIC;�         �      )          rst           : in  STD_LOGIC);�         �      !   component cordic_iter is --{{{�         �            generic(�         �      9             N     : natural := 16; --Ancho de la palabra�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �            port(�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   !   #   �      "          m_valid : out STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   #   %   �      "          m_ready : in  STD_LOGIC;�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   )   +   �      "          s_valid : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   -   /   �      (          clk           : in  STD_LOGIC;�   .   0   �      )          rst           : in  STD_LOGIC);�   /   1   �         end component; --}}}�   1   3   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   2   4   �      8   type   axiStates   is (waitingSvalid, waitingMready);�   3   5   �      1   signal preState  : axiStates := waitingSvalid;�   4   6   �      1   signal posState  : axiStates := waitingSvalid;�   5   7   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   6   8   �      "   signal xyData    : xyDataArray;�   7   9   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   :   <   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   ;   =   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   <   >   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   =   ?   �      A   signal validW, readyW, inv  : handShakeVector:= (others=>'0');�   >   @   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   ?   A   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   B   D   �      )   pre_cordic_proc:process (clk) is --{{{�   C   E   �      1      variable bitCounter :integer range 0 to 8 ;�   D   F   �         begin�   E   G   �            if rising_edge(clk) then�   F   H   �               if rst = '0' then�   G   I   �      +            preState      <= waitingSvalid;�   H   J   �      !            s_axis_tready <= '1';�   I   K   �      !            validW(0)     <= '0';�   J   L   �      !            inv(0)        <= '0';�   K   M   �                  bitCounter    := 0;�   L   N   �               else�   M   O   �                  case preState is�   N   P   �      $               when waitingSvalid =>�   O   Q   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   P   R   �      2                     bitCounter := bitCounter + 1;�   Q   S   �      '                     case bitCounter is�   R   T   �      !                        when 1 =>�   S   U   �      4                          wirex(0) <= (others=>'0');�   T   V   �      5                          if s_axis_tdata(7)='1' then�   U   W   �      -                             inv(0)   <= '1';�   V   X   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   W   Y   �                                else�   X   Z   �      -                             inv(0)   <= '0';�   Y   [   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   Z   \   �      !                          end if;�   [   ]   �      !                        when 2 =>�   \   ^   �      4                          wirey(0) <= (others=>'0');�   ]   _   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   ^   `   �      ,                          if inv(0)='1' then�   _   a   �      8                             if s_axis_tdata(7)='1' then�   `   b   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   a   c   �      "                             else �   b   d   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   c   e   �      $                             end if;�   d   f   �                                else �   e   g   �      7                             wirez(0) <= (others=>'0');�   f   h   �      !                          end if;�   g   i   �      /                          validW(0)     <= '1';�   h   j   �      v                          if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   i   k   �      k                          s_axis_tready <= '0';                           --entonces yo tambien estoy listo�   j   l   �      9                          preState      <= waitingMready;�   k   m   �      &                        when others =>�   l   n   �                           end case;�   m   o   �                        else�   n   p   �      &                     validW(0) <= '0';�   o   q   �                        end if;�   p   r   �      $               when waitingMready =>�   q   s   �      n                  if readyW(0) = '1' then                           --espero e que este listo para enviar algo�   r   t   �      *                     validW(0)     <= '0';�   s   u   �      f                     s_axis_tready <= '1';                           --entonces yo tambien estoy listo�   t   v   �      4                     preState      <= waitingSvalid;�   u   w   �      (                     bitCounter    := 0;�   v   x   �                        end if;�   w   y   �                     when others =>�   x   z   �                  end case;�   y   {   �               end if;�   z   |   �            end if;�   {   }   �      %   end process pre_cordic_proc; --}}}�   }      �      )   pos_cordic_proc:process (clk) is --{{{�   ~   �   �      1      variable bitCounter :integer range 0 to 8 ;�      �   �         begin�   �   �   �            if rising_edge(clk) then�   �   �   �               if rst = '0' then�   �   �   �      +            posState      <= waitingSvalid;�   �   �   �      !            m_axis_tvalid <= '0';�   �   �   �      -            m_axis_tdata  <= (others => '0');�   �   �   �      -            angle         <= (others => '0');�   �   �   �      T            readyW(ITER)  <= '1';                           --y ya no tengo mas nada�   �   �   �                  bitCounter := 0;�   �   �   �               else�   �   �   �                  case posState is�   �   �   �      $               when waitingSvalid =>�   �   �   �      q                  if validW(ITER) = '1' then                           --espero e que este listo para enviar algo�   �   �   �      -                     if(inv(ITER-1)='1') then�   �   �   �      J                        angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      ^                        m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �                           else�   �   �   �      I                        angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �      C                        m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �                           end if;�   �   �   �      *                     readyW(ITER)  <= '0';�   �   �   �      *                     m_axis_tvalid <= '1';�   �   �   �      (                     bitCounter    := 0;�   �   �   �      4                     posState      <= waitingMready;�   �   �   �                        end if;�   �   �   �      '                  when waitingMready =>�   �   �   �      0                     if m_axis_tready = '1' then�   �   �   �      +                        bitCounter    := 0;�   �   �   �      }                        posState      <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      �                        m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      -                        readyW(ITER)  <= '1';�   �   �   �                           end if;�   �   �   �                     end case;�   �   �   �                  end if;�   �   �   �               end if;�   �   �   �      %   end process pos_cordic_proc; --}}}�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �         begin�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �            iteration: cordic_iter�   �   �   �            generic map(N,j)�   �   �   �            port  map (�   �   �   �      '           m_dataX => wirex    ( j+1 ),�   �   �   �      '           m_dataY => wirey    ( j+1 ),�   �   �   �      '           m_dataZ => wirez    ( j+1 ),�   �   �   �      '           m_valid => validW   ( j+1 ),�   �   �   �      '           m_inv   => inv      ( j+1 ),�   �   �   �      '           m_ready => readyW   ( j+1 ),�   �   �   �      '           s_dataX => wirex    ( j   ),�   �   �   �      '           s_dataY => wirey    ( j   ),�   �   �   �      '           s_dataZ => wirez    ( j   ),�   �   �   �      '           s_dataT => wireLUT  ( j   ),�   �   �   �      '           s_valid => validW   ( j   ),�   �   �   �      '           s_ready => readyW   ( j   ),�   �   �   �      '           s_inv   => inv      ( j   ),�   �   �   �                 clk     => clk,�   �   �   �                 rst     => rst�   �   �   �               );�   �   �   �         end generate;5�_�  W  Y      Z  X   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�     �   �   �   �    �   �   �   �                           end if;   *                     readyW(ITER)  := '0';5�_�  X              Y   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�     �   �   �                            end if;5�_�  J          L  K   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^��     �   �   �        5�_�  H          J  I   �       ����                                                                                                                                                                >   
                                                       �                                                                                              �          �          V       ^�`     �   �   �   �                           �   �   �   �      &                     kkkkkkkkkkkkkkkkk5�_�  �  �  �  �  �   y        ����                                                                                                                                                                >   
                                                       �                                                                                              y           y           V        ^�8     �   x   |        5�_�  �              �   y       ����                                                                                                                                                                >   
                                                       �                                                                                              {          |          V       ^�9     �   x   z        5�_�  �          �  �   y        ����                                                                                                                                                                >   
                                                       �                                                                                              y           y          V       ^�5     �   x   ~        5�_�  �      �  �  �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   y   {   �      h                  if ER) = '1' then                           --espero e que este listo para enviar algo5�_�  �          �  �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              z                           ^�     �   y   {   �      m                  if validER) = '1' then                           --espero e que este listo para enviar algo5�_�  �          �  �   z       ����                                                                                                                                                                >   
                                                       �                                                                                              x          y          V       ^��     �   y   {   �      t                  -if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  �          �  �   y   "    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��   �   x   z   �      u                  if m_readyW(ITER-1) = '1' then                           --espero e que este listo para enviar algo5�_�  �          �  �   y   "    ����                                                                                                                                                                                                                            �                                                                                              K           T           V        ^��     �   x   z   �      s                  if m_readyW(ITER) = '1' then                           --espero e que este listo para enviar algo5�_�  &          (  '   T        ����                                                                                                                                                                                                                                                                                                                            �          �   !       V   !    ^q"     �   T   U   �    �   S   T   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada5�_�  �          �  �   �        ����                                                                                                                                                                                                                                                                                                                            �          �          V       ^n�     �   �   �          #      port                     map(�   �   �          2                 m_dataX       => wirex   ( j+1 ),�   �   �          2                 m_dataY       => wirey   ( j+1 ),�   �   �          2                 m_dataZ       => wirez   ( j+1 ),�   �   �          2                 m_valid       => dv      ( j   ),�   �   �          2                 m_inv         => inv     ( j+1 ),�   �   �          !                 m_ready       =>�   �   �          2                    s_dataX    => wirex   ( j   ),�   �   �          2                    s_dataY    => wirey   ( j   ),�   �   �          2                    s_dataZ    => wirez   ( j   ),�   �   �          2                    s_dataT    => wireLUT ( j   ),�   �   �          !                    s_valid    =>�   �   �          2                       s_ready => en      ( j   ),�   �   �          2                       s_inv   => inv     ( j   ),�   �   �          !                       s_atan  =>�   �   �          &                          clk  => clk,�   �   �          %                          rst  => rst�         �         generic(�         �      9             N     : natural := 16; --Ancho de la palabra�      	   �      I             ITER  : natural := 10); -- numero de iteraciones por defecto�      
   �         Port(�   	      �      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);�   
      �      (          m_axis_tvalid : out STD_LOGIC;�         �      (          m_axis_tlast  : out STD_LOGIC;�         �      (          m_axis_tready : in  STD_LOGIC;�         �      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);�         �      (          s_axis_tvalid : in  STD_LOGIC;�         �      (          s_axis_tlast  : in  STD_LOGIC;�         �      (          s_axis_tready : out STD_LOGIC;�         �      (          clk           : in  STD_LOGIC;�         �      )          rst           : in  STD_LOGIC);�         �      !   component cordic_iter is --{{{�         �            generic(�         �      9             N     : natural := 16; --Ancho de la palabra�         �      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         �            port(�          �      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      !   �      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�       "   �      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   !   #   �      "          m_valid : out STD_LOGIC;�   "   $   �      "          m_inv   : out STD_LOGIC;�   #   %   �      "          m_ready : in  STD_LOGIC;�   %   '   �      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�   &   (   �      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�   '   )   �      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�   (   *   �      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�   )   +   �      "          s_valid : in  STD_LOGIC;�   *   ,   �      "          s_ready : out STD_LOGIC;�   +   -   �      "          s_inv   : in  STD_LOGIC;�   ,   .   �      "          s_atan  : in  STD_LOGIC;�   .   0   �      (          clk           : in  STD_LOGIC;�   /   1   �      )          rst           : in  STD_LOGIC);�   0   2   �                );�   1   3   �         end component; --}}}�   3   5   �      d   constant MAX_ITER : natural := 10;  -- maximo largo de la tabla. ITER puede ir de aca para abajo �   4   6   �      F   type   axiStates   is (waitingSvalid, waitingMready,waitingCordic);�   5   7   �      1   signal state     : axiStates := waitingSvalid;�   6   8   �      K   type   xyDataArray is array (0 to 1) of std_logic_vector ( 7 downto 0 );�   7   9   �      "   signal xyData    : xyDataArray;�   8   :   �      '   signal clockWise : std_logic := '0';�   9   ;   �      E   signal angle     : std_logic_vector(N-1 downto 0):= (others=>'0');�   :   <   �         �   <   >   �      V   type   handShakeVector is array ( ITER downto 0 )of std_logic                     ;�   =   ?   �      V   type   ConnectVector is array   ( ITER downto 0 )of std_logic_vector(N-1 downto 0);�   >   @   �      �   type   intLUT is array          ( MAX_ITER-1 downto 0 )of integer range 0 to 5000  ; --la tabla soporta hasta MAX_ITER, pero en la instanciacino del cordic se puede elejir menos o igual.. no mas porque reviente.. la tabla no tendria datos..�   ?   A   �      C   signal en, dv, inv            : handShakeVector:= (others=>'0');�   @   B   �      6   signal wirex, wirey, wirez, wireLUT: ConnectVector;�   A   C   �      j   signal atanLUT                     : intLUT       := (4500, 2657, 1404, 713, 358, 179, 90, 45, 22, 11);�   D   F   �      %   cordic_proc:process (clk) is --{{{�   E   G   �      1      variable bitCounter :integer range 0 to 8 ;�   G   I   �      *      variable sign :signed (15 downto 0);�   H   J   �      9      variable extension :std_logic_vector (15 downto 0);�   I   K   �         begin�   J   L   �            if rising_edge(clk) then�   K   M   �               if rst = '0' then�   L   N   �      +            state         <= waitingSvalid;�   M   O   �      !            s_axis_tready <= '1';�   N   P   �      !            m_axis_tvalid <= '0';�   O   Q   �      -            m_axis_tdata  <= (others => '0');�   P   R   �      !            clockWise     <= '0';�   Q   S   �      -            angle         <= (others => '0');�   R   T   �      T            en(0)         <= '0';                           --y ya no tengo mas nada�   S   U   �      T            inv(0)        <= '0';                           --y ya no tengo mas nada�   T   V   �                  bitCounter    := 0;�   U   W   �               else�   V   X   �                  case state is�   W   Y   �      $               when waitingSvalid =>�   X   Z   �      r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo�   Y   [   �      '                     case bitCounter is�   Z   \   �      !                        when 0 =>�   [   ]   �      4                          wirex(0) <= (others=>'0');�   \   ^   �      5                          if s_axis_tdata(7)='1' then�   ]   _   �      -                             inv(0)   <= '1';�   ^   `   �      k                             wirex(0) <= std_logic_vector(to_signed(to_integer(-signed(s_axis_tdata)),16));�   _   a   �                                else�   `   b   �      -                             inv(0)   <= '0';�   a   c   �      j                             wirex(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   b   d   �      !                          end if;�   c   e   �      !                        when 1 =>�   d   f   �      4                          wirey(0) <= (others=>'0');�   e   g   �      g                          wirey(0) <= std_logic_vector(to_signed(to_integer(signed(s_axis_tdata)),16));�   f   h   �      ,                          if inv(0)='1' then�   g   i   �      8                             if s_axis_tdata(7)='1' then�   h   j   �      _                                wirez(0) <= std_logic_vector(to_signed(18000,wirez(0)'length));�   i   k   �      "                             else �   j   l   �      `                                wirez(0) <= std_logic_vector(to_signed(-18000,wirez(0)'length));�   k   m   �      $                             end if;�   l   n   �                                else �   m   o   �      :                                wirez(0) <= (others=>'0');�   n   p   �      !                          end if;�   o   q   �      i                          en(0)                <= '1';                           --y ya no tengo mas nada�   p   r   �      r                          s_axis_tready        <= '0';                           --entonces yo tambien estoy listo�   q   s   �      i                          m_axis_tvalid        <= '0';                           --y ya no tengo mas nada�   r   t   �      @                          state                <= waitingCordic;�   s   u   �      &                        when others =>�   t   v   �                           end case;�   u   w   �      2                     bitCounter := bitCounter + 1;�   v   x   �                        end if;�   w   y   �      $               when waitingCordic =>�   x   z   �      !                  en ( 0 )<= '0';�   y   {   �      j                  if dv(0) = '1' then                           --espero e que este listo para enviar algo�   z   |   �      @                     m_axis_tdata  <= wirex(ITER-1)(7 downto 0);�   {   }   �      ]                     m_axis_tvalid <= '1';                           --y ya no tengo mas nada�   |   ~   �      4                     state         <= waitingMready;�   }      �      (                     bitCounter    := 0;�   ~   �   �                        end if;�   �   �   �      $               when waitingMready =>�   �   �   �      l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?�   �   �   �      N                    bitCounter := bitCounter+1;                   --incremento�   �   �   �      '                     case bitCounter is�   �   �   �      !                        when 1 =>�   �   �   �      E                           m_axis_tdata <= wirey(ITER-1)(7 downto 0);�   �   �   �      !                        when 2 =>�   �   �   �      3                           if(inv(ITER-1)='1') then�   �   �   �      P                              angle <= std_logic_vector(-signed(wirez(ITER-1)));�   �   �   �      d                              m_axis_tdata <= std_logic_vector(-signed(wirez(ITER-1)(14 downto 7)));�   �   �   �                                 else�   �   �   �      O                              angle <= std_logic_vector(signed(wirez(ITER-1)));�   �   �   �      I                              m_axis_tdata <= wirez(ITER-1)(14 downto 7);�   �   �   �      "                           end if;�   �   �   �      �                           m_axis_tvalid <= '0';                      --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar�   �   �   �      0                           s_axis_tready <= '1';�   �   �   �      .                           bitCounter    := 0;�   �   �   �      �                           state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato�   �   �   �      &                        when others =>�   �   �   �                           end case;�   �   �   �                        end if;�   �   �   �                  end case;�   �   �   �               end if;�   �   �   �            end if;�   �   �   �      !   end process cordic_proc; --}}}�   �   �   �      5   connection_instance: for j in 0 to ITER-1 generate�   �   �   �         begin�   �   �   �      G      wireLUT(j) <= std_logic_vector(to_unsigned(atanLUT(ITER-1-j),N));�   �   �   �            iteration: cordic_iter�   �   �   �            generic map(N,j)�   �   �   �      #      port                     map(�   �   �   �      2                 m_dataX       => wirex   ( j+1 ),�   �   �   �      2                 m_dataY       => wirey   ( j+1 ),�   �   �   �      2                 m_dataZ       => wirez   ( j+1 ),�   �   �   �      2                 m_valid       => dv      ( j   ),�   �   �   �      2                 m_inv         => inv     ( j+1 ),�   �   �   �      !                 m_ready       =>�   �   �   �      2                    s_dataX    => wirex   ( j   ),�   �   �   �      2                    s_dataY    => wirey   ( j   ),�   �   �   �      2                    s_dataZ    => wirez   ( j   ),�   �   �   �      2                    s_dataT    => wireLUT ( j   ),�   �   �   �      !                    s_valid    =>�   �   �   �      2                       s_ready => en      ( j   ),�   �   �   �      2                       s_inv   => inv     ( j   ),�   �   �   �      !                       s_atan  =>�   �   �   �      &                          clk  => clk,�   �   �   �      %                          rst  => rst�   �   �   �                             );�   �   �   �               en(j+1)<=dv(j);�   �   �   �         end generate;5�_�  �          �  �   �       ����                                                                                                                                                                                                                                                                                                                            �          �                 ^m�     �   �   �        �   �   �   �       5��