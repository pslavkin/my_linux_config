Vim�UnDo� �+fR�(��"#�����v ��|w�۶�d   A                                   ^�S    _�                     +       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   *   +          V                     --m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                   2       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   1   2          S                     --bitCounter := bitCounter+1;                     --incremento5�_�                    4       ����                                                                                                                                                                                                                                                                                                                                                             ^��    �   3   4          Y                        --m_axis_tdata(0) <= s_axis_tdata(bitCounter);    --pongo el dato5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             ^�R    �                (architecture Behavioral of split_1to8 is�                end split_1to8;�                entity split_1to8 is5�_�                    2       ����                                                                                                                                                                                                                                                                                                                                                             ^��     �   1   3        5��