Vim�UnDo� .��c5��s
H��wR��7�vٝ��Nȥ   Y           "                 ^��   < _�                             ����                                                                                                                                                                                                                                                                                                                                                  V        ^�     �         =    �         =    �                    Port(     =           m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);   )           m_axis_tvalid : out STD_LOGIC;   )           m_axis_tlast  : out STD_LOGIC;   )           m_axis_tready : in  STD_LOGIC;       =           s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);   )           s_axis_tvalid : in  STD_LOGIC;   )           s_axis_tlast  : in  STD_LOGIC;   )           s_axis_tready : out STD_LOGIC;       )           clk           : in  STD_LOGIC;   *           rst           : in  STD_LOGIC);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V        ^�     �         O      !   component cordic_iter is --{{{5�_�                            ����                                                                                                                                                                                                                                                                                                                                                 V        ^�"     �                entity mapper is --{{{5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V        ^�&     �         N      end mapper; --}}}5�_�                           ����                                                                                                                                                                                                                                                                                                                                                 V        ^�*     �                   end component; --}}}5�_�                            ����                                                                                                                                                                                                                                                                                                                                                   V        ^�4     �                F   type real_im_array is array (0 to 15) of integer range -128 to 127;   �   constant real_table : real_im_array := (125 ,106 ,71  ,25  ,-25 ,-71 ,-106 ,-125 ,-125 ,-106 ,-71  ,-25  ,25   ,71   ,106 ,125);   �   constant im_table   : real_im_array  := (25  ,71  ,106 ,125 ,125 ,106 ,71   ,25   ,-25  ,-71  ,-106 ,-125 ,-125 ,-106 ,-71 ,-25);       4   type axiStates is (waitingSvalid, waitingMready);   2   signal state      : axiStates := waitingSvalid;   7   signal data2Map   :std_logic_vector ( 3 downto 0 ) ;    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  V        ^�8     �         E         mapper_proc:process (clk) is5�_�      	                 
    ����                                                                                                                                                                                                                                                                                                                                                  V        ^�<     �         E         cordic_proc:process (clk) is5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                                                V       ^�A     �                1      variable bitCounter :integer range 0 to 8 ;   1      variable index      :integer range 0 to 15;5�_�   	              
           ����                                                                                                                                                                                                                                                                                                                                       !           V        ^�O     �      "   ?    �         ?    �                +            state         <= waitingSvalid;   !            s_axis_tready <= '1';   !            m_axis_tvalid <= '0';   -            m_axis_tdata  <= (others => '0');5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                      !                 ^�X     �      "   C      9             xip1  : out std_logic_vector (N-1 downto 0);   9             yip1  : out std_logic_vector (N-1 downto 0);   8             zip1  : out std_logic_vector (N-1 downto 0)�         C      #             dv_o  : out std_logic;5�_�                       $    ����                                                                                                                                                                                                                                                                                                                               $       !   J       ���    ^�}     �      "   C      5             dv_o  <= (others=>'0');;: out std_logic;   K             xip1  <= (others=>'0');;: out std_logic_vector (N-1 downto 0);   K             yip1  <= (others=>'0');;: out std_logic_vector (N-1 downto 0);   J             zip1  <= (others=>'0');;: out std_logic_vector (N-1 downto 0)5�_�                    #        ����                                                                                                                                                                                                                                                                                                                            #          #          V   #    ^��     �   "   $   B    �   #   $   B    �   "   #                      case state is5�_�                    $        ����                                                                                                                                                                                                                                                                                                                            $          >          V       ^��     �   #   $          $               when waitingSvalid =>   r                  if s_axis_tvalid = '1' then                           --espero e que este listo para enviar algo   ?                     data2Map(bitCounter)   <= s_axis_tdata(0);   ?                     data2Map(bitCounter+1) <= s_axis_tdata(1);   >                     bitCounter             := bitCounter + 2;   \                     if bitCounter = 4 then                             --porque bit voy?      H                        index         := to_integer(unsigned(data2Map));   Z                        m_axis_tdata  <= std_logic_vector(to_signed(real_table(index),8));   l                        s_axis_tready <= '0';                              --entonces yo tambien estoy listo   `                        m_axis_tvalid <= '1';                           --y ya no tengo mas nada   +                        bitCounter    := 0;   7                        state         <= waitingMready;                        end if;                     end if;   $               when waitingMready =>   l                  if m_axis_tready = '1' then                      --lo puedo empezar a mandar al otro lado?   O                     bitCounter := bitCounter+1;                   --incremento   a                     if bitCounter < 2 then                        --perfecto, porque bit voy?      X                        m_axis_tdata  <= std_logic_vector(to_signed(im_table(index),8));                        else   �                        m_axis_tvalid <= '0' ;                     --y aviso que no tengo mas nada que mandar state         <= waitingSvalid;                 --termine de mandar, vuelvo a esperar   -                        s_axis_tready <= '1';   +                        bitCounter    := 0;   }                        state         <= waitingSvalid;            --cambio de estado, y le doy un clk para que ponga el dato                        end if;                     end if;               end case;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �         (      $             dv_o  <= (others=>'0');5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       ^��    �         (                   dv_o  <= '0');5�_�                    &       ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �   %   '   (         end process mapper_proc;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       ^��    �         (      $architecture Behavioral of mapper is5�_�                    #       ����                                                                                                                                                                                                                                                                                                                                                v       ^��    �   "   $   (      $             zip1  <= (others=>'0');5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�	    �   "   $   (      -             zip1  <= "1010" & (others=>'0');5�_�                    #        ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�    �   "   $   (      $             zip1  <= (others=>'0');5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�0     �   "   $   (      $             zip1  <= (others=>'1');5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�:     �   "   $   (      (            if(enzip1  <= (others=>'1');5�_�                   #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�D     �   "   %   (      -            if(en_i = zip1  <= (others=>'1');5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�N     �   "   $   )                  if(en_i = '1' then5�_�                    #       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�O     �   #   %   *                     �   #   %   )    5�_�                    $       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�^     �   $   &   *    5�_�                           ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�f     �         ,         �         +    5�_�                       6    ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �         ,    5�_�                            ����                                                                                                                                                                                                                                                                                                                            %          %          v       ^��     �         -      7   type state is array of (waitingValid,waitingEnable);5�_�      !                       ����                                                                                                                                                                                                                                                                                                                            %          %          v       ^��     �         -       5�_�       "           !   $       ����                                                                                                                                                                                                                                                                                                                            %          %          v       ^��     �   #   %   -    �   $   %   -    5�_�   !   #           "   $       ����                                                                                                                                                                                                                                                                                                                            &          &          v       ^��     �   #   %   .      .   variable state: stateType := waitingEnable;5�_�   "   $           #   $       ����                                                                                                                                                                                                                                                                                                                            &          &          v       ^��     �   #   %   .      7            variable state: stateType := waitingEnable;5�_�   #   %           $   $   
    ����                                                                                                                                                                                                                                                                                                                            &          &          v       ^��     �   #   %          .            state: stateType := waitingEnable;5�_�   $   '           %   $       ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   #   %   .      /             state: stateType := waitingEnable;5�_�   %   (   &       '   %       ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   %   (   /                  �   %   '   .    5�_�   '   )           (   *        ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   )   +   0       5�_�   (   *           )   '   "    ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   &   )   0      "               when waitinEnable =5�_�   )   +           *   (        ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   '   (           5�_�   *   ,           +   (        ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   (   *                         dv_o <= '1';�   '   )                      if en_i = '1' then5�_�   +   -           ,   )       ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   )   +   1                           �   )   +   0    5�_�   ,   .           -   *   #    ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   )   +   1      )                     state:=waitingValidi5�_�   -   /           .   *   #    ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   )   +   1      #                     state:=waiting5�_�   .   0           /   *   (    ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   )   +   1      (                     state:=waitingValid5�_�   /   1           0   *   (    ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^��     �   *   ,   2                           �   *   ,   1    5�_�   0   2           1   +       ����                                                                                                                                                                                                                                                                                                                            (          )          V       ^�     �   +   -   2    �   +   ,   2    5�_�   1   4           2   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�     �   +   -   3      #               when waitinEnable =>5�_�   2   5   3       4   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�(     �   +   -   3      $               when waitingValid =>5�_�   4   6           5   ,        ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�.     �   ,   .   4                        �   ,   .   3    5�_�   5   7           6   -       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�>     �   -   /   5                        �   -   /   4    5�_�   6   8           7   .   (    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�O     �   .   0   6                        �   .   0   5    5�_�   7   9           8   /       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�T     �   .   /                            ee5�_�   8   :           9   /        ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�U     �   .   /           5�_�   9   ;           :   /       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�U     �   .   /          &               zip1  <= (others=>'1');5�_�   :   <           ;   .   	    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�W     �   .   0   4                        �   .   0   3    5�_�   ;   @           <   '       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�m     �   &   (          #               when waitinEnable =>5�_�   <   A   =       @   -       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��    �   ,   .   4                        dv_o <= '1';5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      ;   type stateType is array of (waitingValid,waitingEnable);5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      :   type stateType is array f (waitingValid,waitingEnable);5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��    �         4      9   type stateType is array  (waitingValid,waitingEnable);5�_�   C   E           D      7    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      8   type stateType is array (waitingValid,waitingEnable);5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      <   type stateType is array (waitingValid,waitingEnable) of ;5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      6   type stateType is (waitingValid,waitingEnable) of ;5�_�   F   H           G      /    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      5   type stateType is waitingValid,waitingEnable) of ;5�_�   G   I           H      /    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��   	 �         4      3   type stateType is waitingValid,waitingEnableof ;5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �         4      0   type stateType is waitingValid,waitingEnable;5�_�   I   K           J      0    ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��   
 �         4      1   type stateType is (waitingValid,waitingEnable;5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��    �         4      .   variable state: stateType := waitingEnable;5�_�   K   M           L   $       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �   #   %   4      $             state := waitingEnable;5�_�   L   N           M   *       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �   )   +   4      )                     state:=waitingValid;5�_�   M   O           N   .       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^��     �   -   /   4      )                  state := waitingEnable;5�_�   N   P           O   -        ����                                                                                                                                                                                                                                                                                                                            -          .          V       ^��     �   1   3   4          end process cordic_iter_proc;�   0   2   4            end if;�   /   1   4               end if;�   .   0   4                  end case;�   -   /   4      )                  state <= waitingEnable;�   ,   .   4                        dv_o  <= '0';�   +   -   4      #               when waitingValid =>�   *   ,   4                        end if;�   )   +   4      )                     state<=waitingValid;�   (   *   4      !                     dv_o <= '1';�   '   )   4      $                  if en_i = '1' then�   &   (   4      $               when waitingEnable =>�   %   '   4                  case state is�   $   &   4               else�   #   %   4      $             state <= waitingEnable;�   "   $   4      $             zip1  <= (others=>'0');�   !   #   4      $             yip1  <= (others=>'0');�       "   4      $             xip1  <= (others=>'0');�      !   4                   dv_o  <= '0';�          4               if rst = '0' then�         4            if rising_edge(clk) then�         4         begin�         4      $   cordic_iter_proc:process (clk) is�         4      ,   signal state: stateType := waitingEnable;�         4      2   type stateType is (waitingValid,waitingEnable);�         4                );�         4      8             zip1  : out std_logic_vector (N-1 downto 0)�         4      9             yip1  : out std_logic_vector (N-1 downto 0);�         4      9             xip1  : out std_logic_vector (N-1 downto 0);�         4      #             dv_o  : out std_logic;�         4      9             ci    : in  std_logic_vector (N-1 downto 0);�         4      9             zi    : in  std_logic_vector (N-1 downto 0);�         4      9             yi    : in  std_logic_vector (N-1 downto 0);�         4      9             xi    : in  std_logic_vector (N-1 downto 0);�         4      #             en_i  : in  std_logic;�   
      4      #             rst   : in  std_logic;�   	      4      #             clk   : in  std_logic;�      
   4            port(�      	   4      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         4      9             N     : natural := 16; --Ancho de la palabra�         4            generic(�   ,   .                            dv_o <= '0';�   -   /          )                  state <= waitingEnable;5�_�   O   Q           P   )        ����                                                                                                                                                                                                                                                                                                                            )           *           V        ^��    �   1   3   4          end process cordic_iter_proc;�   0   2   4            end if;�   /   1   4               end if;�   .   0   4                  end case;�   -   /   4      )                  state <= waitingEnable;�   ,   .   4                        dv_o  <= '0';�   +   -   4      #               when waitingValid =>�   *   ,   4                        end if;�   )   +   4      +                     state <= waitingValid;�   (   *   4      "                     dv_o  <= '1';�   '   )   4      $                  if en_i = '1' then�   &   (   4      $               when waitingEnable =>�   %   '   4                  case state is�   $   &   4               else�   #   %   4      $             state <= waitingEnable;�   "   $   4      $             zip1  <= (others=>'0');�   !   #   4      $             yip1  <= (others=>'0');�       "   4      $             xip1  <= (others=>'0');�      !   4                   dv_o  <= '0';�          4               if rst = '0' then�         4            if rising_edge(clk) then�         4         begin�         4      $   cordic_iter_proc:process (clk) is�         4      ,   signal state: stateType := waitingEnable;�         4      2   type stateType is (waitingValid,waitingEnable);�         4                );�         4      8             zip1  : out std_logic_vector (N-1 downto 0)�         4      9             yip1  : out std_logic_vector (N-1 downto 0);�         4      9             xip1  : out std_logic_vector (N-1 downto 0);�         4      #             dv_o  : out std_logic;�         4      9             ci    : in  std_logic_vector (N-1 downto 0);�         4      9             zi    : in  std_logic_vector (N-1 downto 0);�         4      9             yi    : in  std_logic_vector (N-1 downto 0);�         4      9             xi    : in  std_logic_vector (N-1 downto 0);�         4      #             en_i  : in  std_logic;�   
      4      #             rst   : in  std_logic;�   	      4      #             clk   : in  std_logic;�      
   4            port(�      	   4      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         4      9             N     : natural := 16; --Ancho de la palabra�         4            generic(�   (   *          !                     dv_o <= '1';�   )   +          )                     state<=waitingValid;5�_�   P   R           Q   &        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�    �   &   /   4      $               when waitingEnable =>   $                  if en_i = '1' then   "                     dv_o  <= '1';   +                     state <= waitingValid;                     end if;   #               when waitingValid =>                     dv_o  <= '0';   )                  state <= waitingEnable;�   %   '   4                  case state is5�_�   Q   S           R   /        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�(    �   .   0   4                  end case;5�_�   R   T           S   &        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�8     �   %   '   4      --            case state is5�_�   S   U           T   &        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�9     �   %   '   4      -            case state is5�_�   T   V           U   '        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�:     �   &   (   4      &--               when waitingEnable =>5�_�   U   W           V   '        ����                                                                                                                                                                                                                                                                                                                            &           .                   ^�:     �   &   (   4      %-               when waitingEnable =>5�_�   V   X           W   (        ����                                                                                                                                                                                                                                                                                                                            (           /                 ^�J    �   '   0   4      &--                  if en_i = '1' then   $--                     dv_o  <= '1';   ---                     state <= waitingValid;   --                  end if;   %--               when waitingValid =>   !--                  dv_o  <= '0';   +--                  state <= waitingEnable;   --            end case;5�_�   W   Y           X   )       ����                                                                                                                                                                                                                                                                                                                            (           /                 ^�r     �   (   *   4    �   )   *   4    5�_�   X   Z           Y   )       ����                                                                                                                                                                                                                                                                                                                            (           0                 ^�t     �   (   *   5      8             zip1  : out std_logic_vector (N-1 downto 0)5�_�   Y   [           Z   )       ����                                                                                                                                                                                                                                                                                                                            (           0                 ^�w     �   (   *   5      @                     zip1  : out std_logic_vector (N-1 downto 0)5�_�   Z   \           [   )   .    ����                                                                                                                                                                                                                                                                                                                            (           0                 ^��    �   (   *   5      S                     zip1  <= (others => '1');: out std_logic_vector (N-1 downto 0)5�_�   [   ]           \   (       ����                                                                                                                                                                                                                                                                                                                            (           0                 ^��     �   (   *   6                           �   (   *   5    5�_�   \   ^           ]   )       ����                                                                                                                                                                                                                                                                                                                            (           1                 ^��     �   (   *   6                           if y5�_�   ]   _           ^   )       ����                                                                                                                                                                                                                                                                                                                            (           1                 ^�j     �   (   *   6                           if yi < 0�   )   *   6    5�_�   ^   `           _   )       ����                                                                                                                                                                                                                                                                                                                            (           1                 ^�l     �   (   *   6                           if0 yi < 05�_�   _   a           `   )       ����                                                                                                                                                                                                                                                                                                                            (           1                 ^�m     �   (   +   6                           if yi < 05�_�   `   b           a   *       ����                                                                                                                                                                                                                                                                                                                            (           2                 ^�r    �   )   +   7                              end if5�_�   a   c           b   )       ����                                                                                                                                                                                                                                                                                                                            (           2                 ^��     �   (   *   7      #                     if yi < 0 then5�_�   b   d           c   )   !    ����                                                                                                                                                                                                                                                                                                                            (           2                 ^��    �   (   *   7      *                     if signed(yi < 0 then5�_�   c   e           d   )       ����                                                                                                                                                                                                                                                                                                                            (           2                 ^��     �   (   *   7      +                     if signed(yi) < 0 then�   )   *   7    5�_�   d   f           e   )       ����                                                                                                                                                                                                                                                                                                                            (           2                 ^��     �   (   *   7      ,                     i0f signed(yi) < 0 then5�_�   e   g           f   )       ����                                                                                                                                                                                                                                                                                                                            (           2                 ^��     �   )   +   7    5�_�   f   h           g   *        ����                                                                                                                                                                                                                                                                                                                            (           3                 ^��     �   *   ,   9                              �   *   ,   8    5�_�   g   i           h   +       ����                                                                                                                                                                                                                                                                                                                            (           4                 ^��     �   *   ,   9                              else�   +   ,   9    5�_�   h   j           i   +       ����                                                                                                                                                                                                                                                                                                                            (           4                 ^��     �   *   ,   9                              e0lse5�_�   i   l           j   +       ����                                                                                                                                                                                                                                                                                                                            (           4                 ^��    �   +   -   9    5�_�   j   m   k       l   )        ����                                                                                                                                                                                                                                                                                                                            )           -           V        ^�     �   )   +   ;                              �   )   +   :    5�_�   l   n           m   *       ����                                                                                                                                                                                                                                                                                                                            )           .           V        ^�     �   )   4   ;    �   *   +   ;    5�_�   m   o           n   *        ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   *   ,             pNew.y=p->y+(p->x>>loop);�   )   +             pNew.x=p->x-(p->y>>loop);5�_�   n   p           o   +       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   *   ,   E      4                           pNew.y=p->y+(p->x>>loop);5�_�   o   q           p   +       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   *   ,   E      3                          pNew.y=p->y+(p->x>>loop);5�_�   p   r           q   +       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   *   ,   E      2                         pNew.y=p->y+(p->x>>loop);5�_�   q   s           r   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      1                        pNew.x=p->x-(p->y>>loop);5�_�   r   t           s   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      0                        New.x=p->x-(p->y>>loop);5�_�   s   u           t   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      /                        ew.x=p->x-(p->y>>loop);5�_�   t   v           u   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      .                        w.x=p->x-(p->y>>loop);5�_�   u   w           v   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      -                        .x=p->x-(p->y>>loop);5�_�   v   x           w   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      ,                        x=p->x-(p->y>>loop);5�_�   w   y           x   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      0                        yip1x=p->x-(p->y>>loop);5�_�   x   z           y   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      /                        yip1=p->x-(p->y>>loop);5�_�   y   {           z   *   !    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      3                        yip1=xip1p->x-(p->y>>loop);5�_�   z   |           {   *   !    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      2                        yip1=xip1->x-(p->y>>loop);5�_�   {   }           |   *   !    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      1                        yip1=xip1>x-(p->y>>loop);5�_�   |   ~           }   *   !    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      0                        yip1=xip1x-(p->y>>loop);5�_�   }              ~   *   #    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      /                        yip1=xip1-(p->y>>loop);5�_�   ~   �              *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      /                        yip1=xip1-(p->y>>loop);5�_�      �           �   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      .                        yip1=xp1-(p->y>>loop);5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      -                        yip1=x1-(p->y>>loop);5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      .                        yip1=xi1-(p->y>>loop);5�_�   �   �           �   *        ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      -                        yip1=xi-(p->y>>loop);5�_�   �   �           �   *   "    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      /                        yip1=xi-yi(p->y>>loop);5�_�   �   �           �   *   #    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�&     �   )   +   E      2                        yip1=xi-yi(15(p->y>>loop);5�_�   �   �           �   *        ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�9     �   )   +   E      D                        yip1=xi-yi(14 downto 0) & yi(15(p->y>>loop);5�_�   �   �           �   *   6    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�Y     �   )   +   E      V                        yip1=xi-yi(15) & y1(15) & yi(14 downto 0) & yi(15(p->y>>loop);5�_�   �   �           �   *   A    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�\     �   )   +   E      V                        yip1=xi-yi(15) & y1(15) & yi(13 downto 0) & yi(15(p->y>>loop);5�_�   �   �           �   *   %    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�     �   )   +   E      B                        yip1=xi-yi(15) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   -    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      O                        yip1=xi-yi(15 downto SHIFT) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   -    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      R                        yip1=xi-yi(15 downto 15-SHIFT) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   -    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      S                        yip1=xi-yi(15 downto *15-SHIFT) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   /    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      S                        yip1=xi-yi(15 downto (15-SHIFT) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   6    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^��     �   )   +   E      S                        yip1=xi-yi(15 downto (14-SHIFT) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   ?    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�7     �   )   +   E      T                        yip1=xi-yi(15 downto (14-SHIFT)) & y1(15) & yi(13 downto 0);5�_�   �   �           �   *   S    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�G     �   )   +   E      h                        yip1=xi-yi(15 downto (14-SHIFT)) & y1(13-SHIFT downto SHIFT5) & yi(13 downto 0);5�_�   �   �           �   *   T    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�H     �   )   +   E      g                        yip1=xi-yi(15 downto (14-SHIFT)) & y1(13-SHIFT downto SHIFT) & yi(13 downto 0);5�_�   �   �           �   *   T    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�H     �   )   +   E      T                        yip1=xi-yi(15 downto (14-SHIFT)) & y1(13-SHIFT downto SHIFT)5�_�   �   �           �   *   >    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�K     �   )   +   E      U                        yip1=xi-yi(15 downto (14-SHIFT)) & y1(13-SHIFT downto SHIFT);5�_�   �   �           �   *   G    ����                                                                                                                                                                                                                                                                                                                            *          +          V       ^�M     �   )   +   E      V                        yip1=xi-yi(15 downto (14-SHIFT)) & y1((13-SHIFT downto SHIFT);5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                            +          5           V       ^�V    �   *   +          1                        pNew.y=p->y+(p->x>>loop);      *p=pNew;      return pNew.y>0;   }   int clock(point_t* p,int loop)   {      point_t pNew;      pNew.x=p->x+(p->y>>loop);      pNew.y=p->y-(p->x>>loop);                           P    5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            +          +           V       ^�]     �   )   +   :      W                        yip1=xi-yi(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   *        ����                                                                                                                                                                                                                                                                                                                            *          *          V       ^�a    �   7   9   :          end process cordic_iter_proc;�   6   8   :            end if;�   5   7   :               end if;�   4   6   :                  end case;�   3   5   :      )                  state <= waitingEnable;�   2   4   :                        dv_o  <= '0';�   1   3   :      #               when waitingValid =>�   0   2   :                        end if;�   /   1   :      +                     state <= waitingValid;�   .   0   :      "                     dv_o  <= '1';�   -   /   :      .                     zip1  <= (others => '1');�   ,   .   :                              end if;�   *   ,   :                              else�   )   +   :      Z                        yip1 <= xi-yi(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);�   (   *   :      +                     if signed(yi) < 0 then�   '   )   :      $                  if en_i = '1' then�   &   (   :      $               when waitingEnable =>�   %   '   :                  case state is�   $   &   :               else�   #   %   :      $             state <= waitingEnable;�   "   $   :      $             zip1  <= (others=>'0');�   !   #   :      $             yip1  <= (others=>'0');�       "   :      $             xip1  <= (others=>'0');�      !   :                   dv_o  <= '0';�          :               if rst = '0' then�         :            if rising_edge(clk) then�         :         begin�         :      $   cordic_iter_proc:process (clk) is�         :      ,   signal state: stateType := waitingEnable;�         :      2   type stateType is (waitingValid,waitingEnable);�         :                );�         :      8             zip1  : out std_logic_vector (N-1 downto 0)�         :      9             yip1  : out std_logic_vector (N-1 downto 0);�         :      9             xip1  : out std_logic_vector (N-1 downto 0);�         :      #             dv_o  : out std_logic;�         :      9             ci    : in  std_logic_vector (N-1 downto 0);�         :      9             zi    : in  std_logic_vector (N-1 downto 0);�         :      9             yi    : in  std_logic_vector (N-1 downto 0);�         :      9             xi    : in  std_logic_vector (N-1 downto 0);�         :      #             en_i  : in  std_logic;�   
      :      #             rst   : in  std_logic;�   	      :      #             clk   : in  std_logic;�      
   :            port(�      	   :      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         :      9             N     : natural := 16; --Ancho de la palabra�         :            generic(�   )   +          X                        yip1<=xi-yi(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   *   %    ����                                                                                                                                                                                                                                                                                                                            *          *          V       ^�_    �   )   +   :      Z                        yip1 <= xi-yi(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            *          *          V       ^�u     �         :    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^�w     �         ;    5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�~     �         <    �         <    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            -          -          V       ^�     �                 5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            ,          ,          V       ^�     �                 5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                            +          +          V       ^��     �         ;      ,   signal state: stateType := waitingEnable;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �         ;      /   signal yisstate: stateType := waitingEnable;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       ^��     �         ;      *   signal yis: stateType := waitingEnable;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^��     �         ;      1   signal yis: signed stateType := waitingEnable;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^��     �         ;         signal yis: signed ;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^��     �         ;         variable yis: signed ;5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^��     �         ;    �         ;    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^��     �                &   variable yis: signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   ;    �   &   '   ;    5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      &   variable yis: signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      /            variable yis: signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      &            yis: signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      '            yis : signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      )            yis :=  signed (15 downto 0);5�_�   �   �           �   &   !    ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      7            yis := (others=> '0') signed (15 downto 0);5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�     �   %   '   <      !            yis := (others=> '0')5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                         /       v   /    ^�    �   %   '   <                  yis := 5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                            &          !          V       ^�      �   $   &          $             state <= waitingEnable;�   #   %          $             zip1  <= (others=>'0');�   "   $          $             yip1  <= (others=>'0');�   !   #          $             xip1  <= (others=>'0');�       "                       dv_o  <= '0';5�_�   �   �   �       �   !        ����                                                                                                                                                                                                                                                                                                                            &          !          V       ^�%     �   9   ;   <          end process cordic_iter_proc;�   8   :   <            end if;�   7   9   <               end if;�   6   8   <                  end case;�   5   7   <      )                  state <= waitingEnable;�   4   6   <                        dv_o  <= '0';�   3   5   <      #               when waitingValid =>�   2   4   <                        end if;�   1   3   <      +                     state <= waitingValid;�   0   2   <      "                     dv_o  <= '1';�   /   1   <      .                     zip1  <= (others => '1');�   .   0   <                              end if;�   ,   .   <                              else�   +   -   <      ^                        yip1 <= xi-yi; --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);�   *   ,   <      +                     if signed(yi) < 0 then�   )   +   <      $                  if en_i = '1' then�   (   *   <      $               when waitingEnable =>�   '   )   <                  case state is�   &   (   <               else�   %   '   <                  yis   := 0;�   $   &   <      #            state <= waitingEnable;�   #   %   <      %            zip1  <= (others => '0');�   "   $   <      %            yip1  <= (others => '0');�   !   #   <      %            xip1  <= (others => '0');�       "   <                  dv_o  <= '0';�      !   <               if rst = '0' then�          <            if rising_edge(clk) then�         <         begin�         <      $   cordic_iter_proc:process (clk) is�         <      &   variable yis: signed (15 downto 0);�         <      ,   signal state: stateType := waitingEnable;�         <      2   type stateType is (waitingValid,waitingEnable);�         <                );�         <      8             zip1  : out std_logic_vector (N-1 downto 0)�         <      9             yip1  : out std_logic_vector (N-1 downto 0);�         <      9             xip1  : out std_logic_vector (N-1 downto 0);�         <      #             dv_o  : out std_logic;�         <      9             ci    : in  std_logic_vector (N-1 downto 0);�         <      9             zi    : in  std_logic_vector (N-1 downto 0);�         <      9             yi    : in  std_logic_vector (N-1 downto 0);�         <      9             xi    : in  std_logic_vector (N-1 downto 0);�         <      #             en_i  : in  std_logic;�   
      <      #             rst   : in  std_logic;�   	      <      #             clk   : in  std_logic;�      
   <            port(�      	   <      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         <      9             N     : natural := 16; --Ancho de la palabra�         <            generic(�       "                      dv_o  <= '0';�   %   '                      yis := 0;�   $   &          #            state <= waitingEnable;�   #   %          #            zip1  <= (others=>'0');�   "   $          #            yip1  <= (others=>'0');�   !   #          #            xip1  <= (others=>'0');5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            +          +          v       ^�-     �   *   ,   <      +                     if signed(yi) < 0 then5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            +          +          v       ^�0     �   *   ,   <      $                     if yi) < 0 then5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            +          +          v       ^�3     �   *   ,   <      $                     if yi) < 0 then5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            +          +          v       ^�4     �   *   ,   <      %                     if yis) < 0 then5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            +          +          v       ^�E     �         <    �         <    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�H     �         =      &   variable yis: signed (15 downto 0);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�I     �         =      %   variable is: signed (15 downto 0);5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�L     �   &   (   =    �   '   (   =    5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                            -          -          v       ^�M     �   '   )   >                  yis   := 0;5�_�   �   �           �   .   "    ����                                                                                                                                                                                                                                                                                                                            -          -          v       ^�Q     �   -   /   >      ^                        yip1 <= xi-yi; --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   &    ����                                                                                                                                                                                                                                                                                                                            -          -          v       ^�S    �   -   /   >      _                        yip1 <= xis-yi; --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^�Y     �                &   variable yis: signed (15 downto 0);   &   variable xis: signed (15 downto 0);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^�[     �         <    �         <    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                V       ^�\    �                &   variable xis: signed (15 downto 0);�                &   variable yis: signed (15 downto 0);5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                            '          (                 ^�v     �   '   )   >                  xis   := 0;�   &   (   >                  yis   := 0;5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�    �   '   )   >      !            xis   := (others=>'0;�   &   (   >      !            yis   := (others=>'0;5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            '           (                   ^��     �   -   /   >      `                        yip1 <= xis-yis; --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   8    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^��    �   -   /   >      q                        yip1 <= std_logic_vector(xis-yis; --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   8    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^��     �   -   /   >      r                        yip1 <= std_logic_vector(xis-yis); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   5    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^��     �   -   /   >      s                        yip1 <= std_logic_vector(xis-yis(); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   D    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�     �   -   /   >                              yip1 <= std_logic_vector(xis-shift_right(yis(); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   J    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�     �   -   /   >      �                        yip1 <= std_logic_vector(xis-shift_right(yis,SHIFT(); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .   K    ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�    �   -   /   >      �                        yip1 <= std_logic_vector(xis-shift_right(yis,SHIFT); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�     �   -   /   >    �   .   /   >    5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            '           (                   ^�     �   .   0   ?      �                        yip1 <= std_logic_vector(xis-shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   .        ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�B     �   -   .          �                        yip1 <= std_logic_vector(xis-shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�C     �   .   0   >    �   /   0   >    5�_�   �   �           �   /   4    ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�L     �   .   0   ?      �                        yip1 <= std_logic_vector(xis-shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   /   4    ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�N     �   .   0   ?    �   /   0   ?    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�P     �   /   1   @      �                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            .          .          V       ^�S     �         @    �         @    5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            /          /          V       ^�T     �          A      )      variable xis: signed (15 downto 0);5�_�   �   �           �   /   N    ����                                                                                                                                                                                                                                                                                                                            /   N       1   �       ���    ^��     �   .   2   A      �                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);   �                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);   �                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT)); --(15 downto (14-SHIFT)) & y1((13-SHIFT) downto SHIFT);5�_�   �   �           �   /   M    ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^��     �   .   2   A      N                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));    N                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));    N                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT)); 5�_�   �   �           �   1   M    ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^��     �   0   2   A      M                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   1   N    ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^��     �   0   2   A      O                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));  5�_�   �   �           �   1   M    ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^��     �   0   2   A      N                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT)); 5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^�     �   0   2   A      M                        zip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   -   "    ����                                                                                                                                                                                                                                                                                                                            /   M       1   M          M    ^�#     �   -   /   B                           �   -   /   A    5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                            0   M       2   M          M    ^�7     �   -   /   B                           yis:=yi5�_�   �   �           �   .   #    ����                                                                                                                                                                                                                                                                                                                            0   M       2   M          M    ^�9     �   -   /   B      #                     yis:=signed(yi5�_�   �   �           �   .   $    ����                                                                                                                                                                                                                                                                                                                            0   M       2   M          M    ^�=     �   -   /   B    �   .   /   B    5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                            1   M       3   M          M    ^�?     �   .   0   C      %                     yis:=signed(yi);5�_�   �   �           �   /   !    ����                                                                                                                                                                                                                                                                                                                            1   M       3   M          M    ^�@     �   .   0   C      %                     xis:=signed(yi);5�_�   �   �           �   /   !    ����                                                                                                                                                                                                                                                                                                                            1   M       3   M          M    ^�B     �   .   0   C    �   /   0   C    5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�C     �   /   1   D      %                     xis:=signed(xi);5�_�   �   �           �   0       ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�I     �   /   1   D      %                     sis:=signed(xi);5�_�   �   �           �   0   !    ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�L     �   /   1   D      %                     zis:=signed(xi);5�_�   �   �           �   0   !    ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�P     �   /   1   D      $                     zis:=signed(c);5�_�   �   �           �   0   #    ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�R     �   /   1   D      &                     zis:=signed(zic);5�_�   �   �           �   0   #    ����                                                                                                                                                                                                                                                                                                                            2   M       4   M          M    ^�_     �   /   1   D    �   0   1   D    5�_�   �   �           �   1       ����                                                                                                                                                                                                                                                                                                                            3   M       5   M          M    ^�`     �   0   2   E      %                     zis:=signed(zi);5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            3   M       5   M          M    ^�c     �   0   2   E      $                     ci:=signed(zi);5�_�   �   �           �   1        ����                                                                                                                                                                                                                                                                                                                            3   M       5   M          M    ^�f     �   0   2   E      #                     ci:=signed(i);5�_�   �   �           �   )        ����                                                                                                                                                                                                                                                                                                                            3   M       5   M          M    ^�j     �   (   *   E    �   )   *   E    5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            4   M       6   M          M    ^��     �   )   +   F      #            xis   := (others=>'0');5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            4   M       6   M          M    ^��     �   )   +   F      "            ci   := (others=>'0');5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                            4   M       6   M          M    ^��     �   (   *   F    �   )   *   F    5�_�   �   �           �   *       ����                                                                                                                                                                                                                                                                                                                            5   M       7   M          M    ^��     �   )   +   G      #            xis   := (others=>'0');5�_�   �   �           �   0        ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^��     �   D   F   G          end process cordic_iter_proc;�   C   E   G            end if;�   B   D   G               end if;�   A   C   G                  end case;�   @   B   G      )                  state <= waitingEnable;�   ?   A   G                        dv_o  <= '0';�   >   @   G      #               when waitingValid =>�   =   ?   G                        end if;�   <   >   G      +                     state <= waitingValid;�   ;   =   G      "                     dv_o  <= '1';�   :   <   G      .                     zip1  <= (others => '1');�   9   ;   G                              end if;�   7   9   G                              else�   6   8   G      P                        zip1 <= zisstd_logic_vector(xis+shift_right(yis,SHIFT));�   5   7   G      M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   4   6   G      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   3   5   G      $                     if yis < 0 then�   2   4   G      '                     ci  := signed(ci);�   1   3   G      '                     zis := signed(zi);�   0   2   G      '                     xis := signed(xi);�   /   1   G      '                     yis := signed(yi);�   .   0   G      $                  if en_i = '1' then�   -   /   G      $               when waitingEnable =>�   ,   .   G                  case state is�   +   -   G               else�   *   ,   G      #            ci    := (others=>'0');�   )   +   G      #            zis   := (others=>'0');�   (   *   G      #            xis   := (others=>'0');�   '   )   G      #            yis   := (others=>'0');�   &   (   G      #            state <= waitingEnable;�   %   '   G      %            zip1  <= (others => '0');�   $   &   G      %            yip1  <= (others => '0');�   #   %   G      %            xip1  <= (others => '0');�   "   $   G                  dv_o  <= '0';�   !   #   G               if rst = '0' then�       "   G            if rising_edge(clk) then�      !   G         begin�          G      )      variable zis: signed (15 downto 0);�         G      )      variable xis: signed (15 downto 0);�         G      )      variable yis: signed (15 downto 0);�         G      $   cordic_iter_proc:process (clk) is�         G      ,   signal state: stateType := waitingEnable;�         G      2   type stateType is (waitingValid,waitingEnable);�         G                );�         G      8             zip1  : out std_logic_vector (N-1 downto 0)�         G      9             yip1  : out std_logic_vector (N-1 downto 0);�         G      9             xip1  : out std_logic_vector (N-1 downto 0);�         G      #             dv_o  : out std_logic;�         G      9             ci    : in  std_logic_vector (N-1 downto 0);�         G      9             zi    : in  std_logic_vector (N-1 downto 0);�         G      9             yi    : in  std_logic_vector (N-1 downto 0);�         G      9             xi    : in  std_logic_vector (N-1 downto 0);�         G      #             en_i  : in  std_logic;�   
      G      #             rst   : in  std_logic;�   	      G      #             clk   : in  std_logic;�      
   G            port(�      	   G      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         G      9             N     : natural := 16; --Ancho de la palabra�         G            generic(�   /   1          %                     yis:=signed(yi);�   0   2          %                     xis:=signed(xi);�   2   4          $                     ci:=signed(ci);�   1   3          %                     zis:=signed(zi);5�_�   �   �           �   7        ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�)     �   6   8   G      P                        zip1 <= zisstd_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   7   4    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�1     �   6   8   G      a                        zip1 <= std_logic_vector(zisstd_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   7   4    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�5     �   6   8   G      b                        zip1 <= std_logic_vector(zis+std_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   7   5    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�8     �   6   8   G      b                        zip1 <= std_logic_vector(zis-std_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   7   5    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�:     �   6   8   G      5                        zip1 <= std_logic_vector(zis-5�_�   �   �           �   7   8    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�?    �   6   8   G      8                        zip1 <= std_logic_vector(zis-ci)5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�G     �   *   ,   G      #            ci    := (others=>'0');5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�H     �   *   ,   G      $            cis    := (others=>'0');5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^�J     �          G    �          G    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^�L     �      !   H      )      variable zis: signed (15 downto 0);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^�M     �      !   H      )      variable xis: signed (15 downto 0);5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^�R     �   3   5   H      '                     ci  := signed(ci);5�_�   �   �           �   8   7    ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^�U    �   7   9   H      9                        zip1 <= std_logic_vector(zis-ci);5�_�   �   �           �   :        ����                                                                                                                                                                                                                                                                                                                            6   5       8   5       V   5    ^�m     �   9   =   H    �   :   ;   H    5�_�   �   �           �   :        ����                                                                                                                                                                                                                                                                                                                            :          <          V       ^�o     �   ;   =          :                        zip1 <= std_logic_vector(zis-cis);�   :   <          M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   9   ;          M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�q     �   H   J   K          end process cordic_iter_proc;�   G   I   K            end if;�   F   H   K               end if;�   E   G   K                  end case;�   D   F   K      )                  state <= waitingEnable;�   C   E   K                        dv_o  <= '0';�   B   D   K      #               when waitingValid =>�   A   C   K                        end if;�   @   B   K      +                     state <= waitingValid;�   ?   A   K      "                     dv_o  <= '1';�   >   @   K      .                     zip1  <= (others => '1');�   =   ?   K                              end if;�   ;   =   K      =                           zip1 <= std_logic_vector(zis-cis);�   :   <   K      P                           yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   9   ;   K      P                           xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   8   :   K                              else�   7   9   K      :                        zip1 <= std_logic_vector(zis-cis);�   6   8   K      M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   5   7   K      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   4   6   K      $                     if yis < 0 then�   3   5   K      '                     cis := signed(ci);�   2   4   K      '                     zis := signed(zi);�   1   3   K      '                     xis := signed(xi);�   0   2   K      '                     yis := signed(yi);�   /   1   K      $                  if en_i = '1' then�   .   0   K      $               when waitingEnable =>�   -   /   K                  case state is�   ,   .   K               else�   +   -   K      #            cis   := (others=>'0');�   *   ,   K      #            zis   := (others=>'0');�   )   +   K      #            xis   := (others=>'0');�   (   *   K      #            yis   := (others=>'0');�   '   )   K      #            state <= waitingEnable;�   &   (   K      %            zip1  <= (others => '0');�   %   '   K      %            yip1  <= (others => '0');�   $   &   K      %            xip1  <= (others => '0');�   #   %   K                  dv_o  <= '0';�   "   $   K               if rst = '0' then�   !   #   K            if rising_edge(clk) then�       "   K         begin�      !   K      )      variable cis: signed (15 downto 0);�          K      )      variable zis: signed (15 downto 0);�         K      )      variable xis: signed (15 downto 0);�         K      )      variable yis: signed (15 downto 0);�         K      $   cordic_iter_proc:process (clk) is�         K      ,   signal state: stateType := waitingEnable;�         K      2   type stateType is (waitingValid,waitingEnable);�         K                );�         K      8             zip1  : out std_logic_vector (N-1 downto 0)�         K      9             yip1  : out std_logic_vector (N-1 downto 0);�         K      9             xip1  : out std_logic_vector (N-1 downto 0);�         K      #             dv_o  : out std_logic;�         K      9             ci    : in  std_logic_vector (N-1 downto 0);�         K      9             zi    : in  std_logic_vector (N-1 downto 0);�         K      9             yi    : in  std_logic_vector (N-1 downto 0);�         K      9             xi    : in  std_logic_vector (N-1 downto 0);�         K      #             en_i  : in  std_logic;�   
      K      #             rst   : in  std_logic;�   	      K      #             clk   : in  std_logic;�      
   K            port(�      	   K      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         K      9             N     : natural := 16; --Ancho de la palabra�         K            generic(�   5   7          M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   7   9          :                        zip1 <= std_logic_vector(zis-cis);�   6   8          M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�   �   �           �   =        ����                                                                                                                                                                                                                                                                                                                            6           8           V        ^�v     �   <   =           5�_�   �              �   :       ����                                                                                                                                                                                                                                                                                                                            :          <                 ^��     �   9   =   J      P                           xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));   P                           yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));   =                           zip1 <= std_logic_vector(zis-cis);5�_�   �                :        ����                                                                                                                                                                                                                                                                                                                            :          <          V       ^��     �   ;   =          :                        zip1 <= std_logic_vector(zis-cis);�   :   <          M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   9   ;          M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));5�_�                  6        ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��   ! �   G   I   J          end process cordic_iter_proc;�   F   H   J            end if;�   E   G   J               end if;�   D   F   J                  end case;�   C   E   J      )                  state <= waitingEnable;�   B   D   J                        dv_o  <= '0';�   A   C   J      #               when waitingValid =>�   @   B   J                        end if;�   ?   A   J      +                     state <= waitingValid;�   >   @   J      "                     dv_o  <= '1';�   =   ?   J      .                     zip1  <= (others => '1');�   <   >   J                              end if;�   ;   =   J      =                           zip1 <= std_logic_vector(zis-cis);�   :   <   J      P                           yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   9   ;   J      P                           xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   8   :   J                              else�   7   9   J      :                        zip1 <= std_logic_vector(zis-cis);�   6   8   J      M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   5   7   J      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   4   6   J      $                     if yis < 0 then�   3   5   J      '                     cis := signed(ci);�   2   4   J      '                     zis := signed(zi);�   1   3   J      '                     xis := signed(xi);�   0   2   J      '                     yis := signed(yi);�   /   1   J      $                  if en_i = '1' then�   .   0   J      $               when waitingEnable =>�   -   /   J                  case state is�   ,   .   J               else�   +   -   J      #            cis   := (others=>'0');�   *   ,   J      #            zis   := (others=>'0');�   )   +   J      #            xis   := (others=>'0');�   (   *   J      #            yis   := (others=>'0');�   '   )   J      #            state <= waitingEnable;�   &   (   J      %            zip1  <= (others => '0');�   %   '   J      %            yip1  <= (others => '0');�   $   &   J      %            xip1  <= (others => '0');�   #   %   J                  dv_o  <= '0';�   "   $   J               if rst = '0' then�   !   #   J            if rising_edge(clk) then�       "   J         begin�      !   J      )      variable cis: signed (15 downto 0);�          J      )      variable zis: signed (15 downto 0);�         J      )      variable xis: signed (15 downto 0);�         J      )      variable yis: signed (15 downto 0);�         J      $   cordic_iter_proc:process (clk) is�         J      ,   signal state: stateType := waitingEnable;�         J      2   type stateType is (waitingValid,waitingEnable);�         J                );�         J      8             zip1  : out std_logic_vector (N-1 downto 0)�         J      9             yip1  : out std_logic_vector (N-1 downto 0);�         J      9             xip1  : out std_logic_vector (N-1 downto 0);�         J      #             dv_o  : out std_logic;�         J      9             ci    : in  std_logic_vector (N-1 downto 0);�         J      9             zi    : in  std_logic_vector (N-1 downto 0);�         J      9             yi    : in  std_logic_vector (N-1 downto 0);�         J      9             xi    : in  std_logic_vector (N-1 downto 0);�         J      #             en_i  : in  std_logic;�   
      J      #             rst   : in  std_logic;�   	      J      #             clk   : in  std_logic;�      
   J            port(�      	   J      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         J      9             N     : natural := 16; --Ancho de la palabra�         J            generic(�   5   7          M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   7   9          :                        zip1 <= std_logic_vector(zis-cis);�   6   8          M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�                 :   =    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�U     �   9   ;   J      P                           xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));5�_�                 ;   4    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�c     �   :   <   J      P                           yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�                 ;   D    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�f     �   :   <   J      P                           yip1 <= std_logic_vector(yis+shift_right(yis,SHIFT));5�_�                 <   7    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�h     �   ;   =   J      =                           zip1 <= std_logic_vector(zis-cis);5�_�                 :   7    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^�}     �   9   ;   J      P                           xip1 <= std_logic_vector(xis-shift+right(yis,SHIFT));5�_�                 ;   7    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��     �   :   <   J      P                           yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));5�_�    	             7   1    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��     �   6   8   J      M                        yip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));5�_�    
          	   7   A    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��     �   6   8   J      M                        yip1 <= std_logic_vector(yis+shift_right(yis,SHIFT));5�_�  	            
   >       ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��   " �   =   >          .                     zip1  <= (others => '1');5�_�  
               :   =    ����                                                                                                                                                                                                                                                                                                                            8          6          V       ^��   # �   9   ;   I      P                           xip1 <= std_logic_vector(xis+shift+right(yis,SHIFT));5�_�                 (        ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��     �   '   (          #            state <= waitingEnable;5�_�                 %       ����                                                                                                                                                                                                                                                                                                                            (          (          V       ^��   ( �   $   &   H    �   %   &   H    5�_�                      ����                                                                                                                                                                                                                                                                                                                                                             ^;x     �         I    �         I    5�_�                        ����                                                                                                                                                                                                                                                                                                                                                       ^;|     �         K      #                 inv_o => inv(j+1),�         K      !                 inv_i => inv(j),5�_�                    &    ����                                                                                                                                                                                                                                                                                                                               &          3       ���    ^;�     �         K      1                 inv_i : in std_logic;l=> inv(j),   3                 inv_o : in std_logic;l=> inv(j+1),5�_�                        ����                                                                                                                                                                                                                                                                                                                               &          3       ���    ^;�     �         K      &                 inv_o : in std_logic;5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       ^;�     �                '                 inv_o : out std_logic;�                &                 inv_i : in std_logic;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                V       ^;�     �         K      "             inv_i : in std_logic;5�_�                         ����                                                                                                                                                                                                                                                                                                                                                V       ^;�     �                #             inv_o : out std_logic;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                V       ^;�   ) �         J    �         J    5�_�                         ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �                #             inv_o : out std_logic;5�_�                        ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�   * �         J    �         J    5�_�                 H        ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �   H   J   L            �   H   J   K    5�_�                 I       ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �   H   J   L            inv_o <5�_�                 I       ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �   H   I                inv_o <=5�_�                 @       ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �   ?   A   K    �   @   A   K    5�_�                 A       ����                                                                                                                                                                                                                                                                                                                                                  V        ^;�     �   @   B   L      "                     dv_o  <= '1';5�_�                  A       ����                                                                                                                                                                                                                                                                                                                            A          A   !       v   !    ^;�     �   @   B   L      #                     inv_o  <= '1';5�_�    !              @        ����                                                                                                                                                                                                                                                                                                                            @   !       B   $       V   $    ^<   + �   I   K   L          end process cordic_iter_proc;�   H   J   L            end if;�   G   I   L               end if;�   F   H   L                  end case;�   E   G   L      )                  state <= waitingEnable;�   D   F   L                        dv_o  <= '0';�   C   E   L      #               when waitingValid =>�   B   D   L                        end if;�   A   C   L      +                     state <= waitingValid;�   @   B   L      %                     inv_o <= inv_in;�   ?   A   L      "                     dv_o  <= '1';�   >   @   L                              end if;�   =   ?   L      =                           zip1 <= std_logic_vector(zis+cis);�   <   >   L      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   ;   =   L      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   :   <   L                              else�   9   ;   L      :                        zip1 <= std_logic_vector(zis-cis);�   8   :   L      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   7   9   L      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   6   8   L      $                     if yis < 0 then�   5   7   L      '                     cis := signed(ci);�   4   6   L      '                     zis := signed(zi);�   3   5   L      '                     xis := signed(xi);�   2   4   L      '                     yis := signed(yi);�   1   3   L      $                  if en_i = '1' then�   0   2   L      $               when waitingEnable =>�   /   1   L                  case state is�   .   0   L               else�   -   /   L      #            cis   := (others=>'0');�   ,   .   L      #            zis   := (others=>'0');�   +   -   L      #            xis   := (others=>'0');�   *   ,   L      #            yis   := (others=>'0');�   )   +   L      %            zip1  <= (others => '0');�   (   *   L      %            yip1  <= (others => '0');�   '   )   L      %            xip1  <= (others => '0');�   &   (   L      #            state <= waitingEnable;�   %   '   L                  dv_o  <= '0';�   $   &   L               if rst = '0' then�   #   %   L            if rising_edge(clk) then�   "   $   L         begin�   !   #   L      )      variable cis: signed (15 downto 0);�       "   L      )      variable zis: signed (15 downto 0);�      !   L      )      variable xis: signed (15 downto 0);�          L      )      variable yis: signed (15 downto 0);�         L      $   cordic_iter_proc:process (clk) is�         L      ,   signal state: stateType := waitingEnable;�         L      2   type stateType is (waitingValid,waitingEnable);�         L                );�         L      8             zip1  : out std_logic_vector (N-1 downto 0)�         L      9             yip1  : out std_logic_vector (N-1 downto 0);�         L      9             xip1  : out std_logic_vector (N-1 downto 0);�         L      #             inv_o : out std_logic;�         L      #             dv_o  : out std_logic;�         L      9             ci    : in  std_logic_vector (N-1 downto 0);�         L      9             zi    : in  std_logic_vector (N-1 downto 0);�         L      9             yi    : in  std_logic_vector (N-1 downto 0);�         L      9             xi    : in  std_logic_vector (N-1 downto 0);�         L      #             inv_i : in  std_logic;�         L      #             en_i  : in  std_logic;�   
      L      #             rst   : in  std_logic;�   	      L      #             clk   : in  std_logic;�      
   L            port(�      	   L      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         L      9             N     : natural := 16; --Ancho de la palabra�         L            generic(�   ?   A          "                     dv_o  <= '1';�   A   C          +                     state <= waitingValid;�   @   B          &                     inv_o  <= inv_in;5�_�     "          !   A   #    ����                                                                                                                                                                                                                                                                                                                            @   !       B   $       V   $    ^<X   - �   @   B   L      %                     inv_o <= inv_in;5�_�  !  #          "   &        ����                                                                                                                                                                                                                                                                                                                            @   !       B   $       V   $    ^>�     �   %   '   L    5�_�  "  $          #   (       ����                                                                                                                                                                                                                                                                                                                            A   !       C   $       V   $    ^>�     �   '   )   M    �   (   )   M    5�_�  #  %          $   (       ����                                                                                                                                                                                                                                                                                                                            B   !       D   $       V   $    ^>�     �   '   )   N                  dv_o  <= '0';5�_�  $  &          %   (       ����                                                                                                                                                                                                                                                                                                                            B   !       D   $       V   $    ^>�     �   '   )   N                  inv_o  <= '0';5�_�  %  '          &   &        ����                                                                                                                                                                                                                                                                                                                            B   !       D   $       V   $    ^>�   . �   %   &           5�_�  &  (          '   )        ����                                                                                                                                                                                                                                                                                                                            /           )           V        ^]_   / �   J   L   M          end process cordic_iter_proc;�   I   K   M            end if;�   H   J   M               end if;�   G   I   M                  end case;�   F   H   M      )                  state <= waitingEnable;�   E   G   M                        dv_o  <= '0';�   D   F   M      #               when waitingValid =>�   C   E   M                        end if;�   B   D   M      +                     state <= waitingValid;�   A   C   M      $                     inv_o <= inv_i;�   @   B   M      "                     dv_o  <= '1';�   ?   A   M                              end if;�   >   @   M      =                           zip1 <= std_logic_vector(zis+cis);�   =   ?   M      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   <   >   M      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   ;   =   M                              else�   :   <   M      :                        zip1 <= std_logic_vector(zis-cis);�   9   ;   M      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   8   :   M      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   7   9   M      $                     if yis < 0 then�   6   8   M      '                     cis := signed(ci);�   5   7   M      '                     zis := signed(zi);�   4   6   M      '                     xis := signed(xi);�   3   5   M      '                     yis := signed(yi);�   2   4   M      $                  if en_i = '1' then�   1   3   M      $               when waitingEnable =>�   0   2   M                  case state is�   /   1   M               else�   .   0   M      $            cis  := (others => '0');�   -   /   M      $            zis  := (others => '0');�   ,   .   M      $            xis  := (others => '0');�   +   -   M      $            yis  := (others => '0');�   *   ,   M      $            zip1 <= (others => '0');�   )   +   M      $            yip1 <= (others => '0');�   (   *   M      $            xip1 <= (others => '0');�   '   )   M      #            state <= waitingEnable;�   &   (   M                  inv_o <= '0';�   %   '   M                  dv_o  <= '0';�   $   &   M               if rst = '0' then�   #   %   M            if rising_edge(clk) then�   "   $   M         begin�   !   #   M      )      variable cis: signed (15 downto 0);�       "   M      )      variable zis: signed (15 downto 0);�      !   M      )      variable xis: signed (15 downto 0);�          M      )      variable yis: signed (15 downto 0);�         M      $   cordic_iter_proc:process (clk) is�         M      ,   signal state: stateType := waitingEnable;�         M      2   type stateType is (waitingValid,waitingEnable);�         M                );�         M      8             zip1  : out std_logic_vector (N-1 downto 0)�         M      9             yip1  : out std_logic_vector (N-1 downto 0);�         M      9             xip1  : out std_logic_vector (N-1 downto 0);�         M      #             inv_o : out std_logic;�         M      #             dv_o  : out std_logic;�         M      9             ci    : in  std_logic_vector (N-1 downto 0);�         M      9             zi    : in  std_logic_vector (N-1 downto 0);�         M      9             yi    : in  std_logic_vector (N-1 downto 0);�         M      9             xi    : in  std_logic_vector (N-1 downto 0);�         M      #             inv_i : in  std_logic;�         M      #             en_i  : in  std_logic;�   
      M      #             rst   : in  std_logic;�   	      M      #             clk   : in  std_logic;�      
   M            port(�      	   M      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         M      9             N     : natural := 16; --Ancho de la palabra�         M            generic(�   (   *          %            xip1  <= (others => '0');�   .   0          #            cis   := (others=>'0');�   -   /          #            zis   := (others=>'0');�   ,   .          #            xis   := (others=>'0');�   +   -          #            yis   := (others=>'0');�   *   ,          %            zip1  <= (others => '0');�   )   +          %            yip1  <= (others => '0');5�_�  '  )          (   
        ����                                                                                                                                                                                                                                                                                                                            /           )           V        ^j     �   	      M    �   
      M    5�_�  (  *          )   
       ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jP     �   	      Y      <          m_axis_tdata  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  )  +          *   
       ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jQ     �   	      Y      =          m_axis_tdatax  : out STD_LOGIC_VECTOR (7 downto 0);5�_�  *  ,          +   
       ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jR     �   	      Y      <          m_axis_tdatax : out STD_LOGIC_VECTOR (7 downto 0);5�_�  +  -          ,          ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^j_     �         Y      <          s_axis_tdata  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  ,  .          -          ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^j_     �         Y      =          s_axis_tdataX  : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  -  /          .      0    ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jc     �         Y      <          s_axis_tdataX : in  STD_LOGIC_VECTOR (7 downto 0);5�_�  .  0          /      3    ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^je     �         Y      ?          s_axis_tdataX : in  STD_LOGIC_VECTOR (N-17 downto 0);5�_�  /  1          0   
   0    ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jh     �   	      Y      <          m_axis_tdataX : out STD_LOGIC_VECTOR (7 downto 0);5�_�  0  2          1   
   3    ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jj     �   	      Y      ?          m_axis_tdataX : out STD_LOGIC_VECTOR (N-17 downto 0);5�_�  1  3          2   
       ����                                                                                                                                                                                                                                                                                                                            ;           5           V        ^jl     �   	      Y    �   
      Y    5�_�  2  4          3   
   
    ����                                                                                                                                                                                                                                                                                                                            <           6           V        ^jl     �   	      Z    �   
      Z    5�_�  3  5          4          ����                                                                                                                                                                                                                                                                                                                            =           7           V        ^jo     �   
      [      >          m_axis_tdataX : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  4  6          5          ����                                                                                                                                                                                                                                                                                                                            =           7           V        ^jp     �         [      >          m_axis_tdataX : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  5  7          6          ����                                                                                                                                                                                                                                                                                                                            =           7           V        ^jv     �         [    �         [    5�_�  6  8          7          ����                                                                                                                                                                                                                                                                                                                            >           8           V        ^jw     �         \    �         \    5�_�  7  9          8          ����                                                                                                                                                                                                                                                                                                                            ?           9           V        ^jz     �         ]      >          s_axis_tdataX : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  8  :          9          ����                                                                                                                                                                                                                                                                                                                            ?           9           V        ^j|     �         ]      >          s_axis_tdataX : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  9  ;          :          ����                                                                                                                                                                                                                                                                                                                            ?           9           V        ^j     �         ]      >          m_axis_tdataz : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  :  <          ;           ����                                                                                                                                                                                                                                                                                                                            ?           9           V        ^j�     �         ]    �         ]    5�_�  ;  =          <          ����                                                                                                                                                                                                                                                                                                                            @           :           V        ^j�     �         ^      (          s_axis_tlast  : in  STD_LOGIC;5�_�  <  >          =          ����                                                                                                                                                                                                                                                                                                                            @           :           V        ^j�     �         ^      (          s_axis_tquad  : in  STD_LOGIC;5�_�  =  ?          >          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      >          s_axis_tdataY : in  STD_LOGIC_VECTOR (N-1 downto 0);   >          s_axis_tdataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);   (          s_axis_tvalid : in  STD_LOGIC;   (          s_axis_tlast  : in  STD_LOGIC;   (          s_axis_tready : out STD_LOGIC;�         ^      >          s_axis_tdataX : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  >  @          ?          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      -          s_axis_tcuadrante  : in  STD_LOGIC;5�_�  ?  A          @          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      .          s_axis_tcuadrante   : in  STD_LOGIC;5�_�  @  B          A          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      *          s_axis_tinver   : in  STD_LOGIC;5�_�  A  C          B          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      )          s_axis_tinver  : in  STD_LOGIC;5�_�  B  D          C          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      D          s_axis_tdataX       : in  STD_LOGIC_VECTOR (N-1 downto 0);   D          s_axis_tdataY       : in  STD_LOGIC_VECTOR (N-1 downto 0);   D          s_axis_tdataZ       : in  STD_LOGIC_VECTOR (N-1 downto 0);   .          s_axis_tvalid       : in  STD_LOGIC;   .          s_axis_tlast        : in  STD_LOGIC;   .          s_axis_tready       : out STD_LOGIC;5�_�  C  E          D          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      C          s_axis_tdataX      : in  STD_LOGIC_VECTOR (N-1 downto 0);   C          s_axis_tdataY      : in  STD_LOGIC_VECTOR (N-1 downto 0);   C          s_axis_tdataZ      : in  STD_LOGIC_VECTOR (N-1 downto 0);   -          s_axis_tvalid      : in  STD_LOGIC;   -          s_axis_tlast       : in  STD_LOGIC;   -          s_axis_tready      : out STD_LOGIC;5�_�  D  F          E          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      (          s_axis_tinver : in  STD_LOGIC;5�_�  E  G          F          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      '          s_axis_tinvr : in  STD_LOGIC;5�_�  F  H          G          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^      &          s_axis_tinv : in  STD_LOGIC;5�_�  G  I          H           ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         ^    �         ^    5�_�  H  J          I          ����                                                                                                                                                                                                                                                                                                                                                       ^j�     �         _      (          s_axis_tinv   : in  STD_LOGIC;5�_�  I  K          J           ����                                                                                                                                                                                                                                                                                                                                                V       ^j�     �                )          s_axis_tinv   : out  STD_LOGIC;5�_�  J  L          K           ����                                                                                                                                                                                                                                                                                                                                                V       ^j�     �         ^    �         ^    5�_�  K  M          L          ����                                                                                                                                                                                                                                                                                                                                                V       ^j�     �         _      )          s_axis_tinv   : out  STD_LOGIC;5�_�  L  N          M           ����                                                                                                                                                                                                                                                                                                                                       (                   ^j�     �      )   _      #             rst   : in  std_logic;   #             en_i  : in  std_logic;   #             inv_i : in  std_logic;   9             xi    : in  std_logic_vector (N-1 downto 0);   9             yi    : in  std_logic_vector (N-1 downto 0);   9             zi    : in  std_logic_vector (N-1 downto 0);   9             ci    : in  std_logic_vector (N-1 downto 0);   #             dv_o  : out std_logic;   #             inv_o : out std_logic;   9             xip1  : out std_logic_vector (N-1 downto 0);   9             yip1  : out std_logic_vector (N-1 downto 0);   8             zip1  : out std_logic_vector (N-1 downto 0)�         _      #             clk   : in  std_logic;5�_�  M  O          N      
    ����                                                                                                                                                                                                                                                                                                                            
                           ^k     �         _      (          s_axis_tinv   : out STD_LOGIC;5�_�  N  P          O   
       ����                                                                                                                                                                                                                                                                                                                            
                           ^k      �   	      _      >          m_axis_tdataX : out STD_LOGIC_VECTOR (N-1 downto 0);   >          m_axis_tdataY : out STD_LOGIC_VECTOR (N-1 downto 0);   >          m_axis_tdataZ : out STD_LOGIC_VECTOR (N-1 downto 0);   (          m_axis_tvalid : out STD_LOGIC;   (          m_axis_tlast  : out STD_LOGIC;   (          m_axis_tinv   : out STD_LOGIC;   (          m_axis_tready : in  STD_LOGIC;5�_�  O  Q          P   
       ����                                                                                                                                                                                                                                                                                                                            
                           ^k"     �   	      _      9          m_tdataX : out STD_LOGIC_VECTOR (N-1 downto 0);   9          m_tdataY : out STD_LOGIC_VECTOR (N-1 downto 0);   9          m_tdataZ : out STD_LOGIC_VECTOR (N-1 downto 0);   #          m_tvalid : out STD_LOGIC;   #          m_tlast  : out STD_LOGIC;   #          m_tinv   : out STD_LOGIC;   #          m_tready : in  STD_LOGIC;5�_�  P  R          Q      
    ����                                                                                                                                                                                                                                                                                                                            
                           ^k$     �                "          m_last  : out STD_LOGIC;5�_�  Q  S          R          ����                                                                                                                                                                                                                                                                                                                                                       ^k)     �         ^      >          s_axis_tdataX : in  STD_LOGIC_VECTOR (N-1 downto 0);   >          s_axis_tdataY : in  STD_LOGIC_VECTOR (N-1 downto 0);   >          s_axis_tdataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);   (          s_axis_tvalid : in  STD_LOGIC;   (          s_axis_tlast  : in  STD_LOGIC;   (          s_axis_tready : out STD_LOGIC;   (          s_axis_tinv   : in  STD_LOGIC;5�_�  R  T          S          ����                                                                                                                                                                                                                                                                                                                                                       ^k+     �         ^      9          s_tdataX : in  STD_LOGIC_VECTOR (N-1 downto 0);   9          s_tdataY : in  STD_LOGIC_VECTOR (N-1 downto 0);   9          s_tdataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);   #          s_tvalid : in  STD_LOGIC;   #          s_tlast  : in  STD_LOGIC;   #          s_tready : out STD_LOGIC;   #          s_tinv   : in  STD_LOGIC;5�_�  S  U          T      
    ����                                                                                                                                                                                                                                                                                                                                                       ^k-     �                "          s_last  : in  STD_LOGIC;5�_�  T  V          U   +       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^k7     �   *   ,   ]      2   type stateType is (waitingValid,waitingEnable);5�_�  U  W          V   ,       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^k:     �   +   -   ]      ,   signal state: stateType := waitingEnable;5�_�  V  X          W   /       ����                                                                                                                                                                                                                                                                                                                            /          2                 ^kJ     �   .   3   ]      )      variable yis: signed (15 downto 0);   )      variable xis: signed (15 downto 0);   )      variable zis: signed (15 downto 0);   )      variable cis: signed (15 downto 0);5�_�  W  Y          X          ����                                                                                                                                                                                                                                                                                                                            /          2                 ^kb     �         ]    �         ]    5�_�  X  Z          Y          ����                                                                                                                                                                                                                                                                                                                            0          3                 ^kc     �         ^      "          s_inv   : in  STD_LOGIC;5�_�  Y  [          Z          ����                                                                                                                                                                                                                                                                                                                            0          3                 ^ke     �         ^      #          s_atan   : in  STD_LOGIC;5�_�  Z  \          [          ����                                                                                                                                                                                                                                                                                                                            0          3                 ^ke     �         ^      "          s_atan  : in  STD_LOGIC;5�_�  [  ]          \          ����                                                                                                                                                                                                                                                                                                                            0          3                 ^kg     �         ^      !          s_atan : in  STD_LOGIC;5�_�  \  ^          ]   3       ����                                                                                                                                                                                                                                                                                                                            0          3                 ^kp     �   2   4   ^      )      variable c_s: signed (15 downto 0);5�_�  ]  _          ^   3       ����                                                                                                                                                                                                                                                                                                                            0          3                 ^kq     �   2   4   ^      -      variable atanc_s: signed (15 downto 0);5�_�  ^  `          _   0       ����                                                                                                                                                                                                                                                                                                                            0          2                 ^kt     �   0   3   ^      )      variable x_s: signed (15 downto 0);   )      variable z_s: signed (15 downto 0);�   /   1   ^      )      variable y_s: signed (15 downto 0);5�_�  _  a          `   3       ����                                                                                                                                                                                                                                                                                                                            0          2                 ^kx     �   2   4   ^      ,      variable atan_s: signed (15 downto 0);5�_�  `  b          a   0       ����                                                                                                                                                                                                                                                                                                                            2          0                 ^k|     �   0   3   ^      .      variable x_signed: signed (15 downto 0);   .      variable z_signed: signed (15 downto 0);�   /   1   ^      .      variable y_signed: signed (15 downto 0);5�_�  a  c          b   3       ����                                                                                                                                                                                                                                                                                                                            2          0                 ^k~     �   2   4   ^      1      variable atan_signed: signed (15 downto 0);5�_�  b  d          c   0   %    ����                                                                                                                                                                                                                                                                                                                            0   %       3   %          %    ^k�     �   0   4   ^      2      variable x_signed    : signed (15 downto 0);   2      variable z_signed    : signed (15 downto 0);   2      variable atan_signed : signed (15 downto 0);�   /   1   ^      2      variable y_signed    : signed (15 downto 0);5�_�  c  f          d   0   (    ����                                                                                                                                                                                                                                                                                                                            0   (       3   )          )    ^k�     �   /   4   ^      5      variable y_signed    : signed (N-115 downto 0);   5      variable x_signed    : signed (N-115 downto 0);   5      variable z_signed    : signed (N-115 downto 0);   5      variable atan_signed : signed (N-115 downto 0);5�_�  d  g  e      f   7       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   6   8   ^                  dv_o  <= '0';5�_�  f  h          g   8       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   7   9   ^                  inv_o <= '0';5�_�  g  i          h   8       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   7   9   ^                  s_inv_o <= '0';5�_�  h  j          i   8       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   7   9   ^                  s_invo <= '0';5�_�  i  k          j   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      $            xip1 <= (others => '0');5�_�  j  l          k   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      '            m_Xxip1 <= (others => '0');5�_�  k  m          l   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      +            m_dataXxip1 <= (others => '0');5�_�  l  n          m   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      *            m_dataXip1 <= (others => '0');5�_�  m  o          n   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      )            m_dataXp1 <= (others => '0');5�_�  n  p          o   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^      (            m_dataX1 <= (others => '0');5�_�  o  q          p   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   ^    �   :   ;   ^    5�_�  p  r          q   :       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   9   ;   _    �   :   ;   _    5�_�  q  s          r   ;       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   :   <   `      '            m_dataX <= (others => '0');5�_�  r  t          s   <       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   ;   =   `      '            m_dataX <= (others => '0');5�_�  s  u          t   <       ����                                                                                                                                                                                                                                                                                                                               
                 v       ^k�     �   ;   =   `      '            m_dataA <= (others => '0');5�_�  t  v          u   =        ����                                                                                                                                                                                                                                                                                                                            =          >          V       ^k�     �   <   =          $            yip1 <= (others => '0');   $            zip1 <= (others => '0');5�_�  u  w          v   =       ����                                                                                                                                                                                                                                                                                                                            =          @                 ^k�     �   =   A   ^      $            xis  := (others => '0');   $            zis  := (others => '0');   $            cis  := (others => '0');�   <   >   ^      $            yis  := (others => '0');5�_�  v  x          w   @       ����                                                                                                                                                                                                                                                                                                                            =          @                 ^k�     �   ?   A   ^      +            c_signedis  := (others => '0');5�_�  w  y          x   @       ����                                                                                                                                                                                                                                                                                                                            =          @                 ^k�     �   ?   A   ^      /            atanc_signedis  := (others => '0');5�_�  x  z          y   @       ����                                                                                                                                                                                                                                                                                                                            =          @                 ^k�     �   ?   A   ^      .            atan_signedis  := (others => '0');5�_�  y  {          z   @       ����                                                                                                                                                                                                                                                                                                                            =          @                 ^k�     �   ?   A   ^      -            atan_signeds  := (others => '0');5�_�  z  |          {   =       ����                                                                                                                                                                                                                                                                                                                            ?          =                 ^k�     �   <   @   ^      +            y_signedis  := (others => '0');   +            x_signedis  := (others => '0');   +            z_signedis  := (others => '0');5�_�  {  }          |   =       ����                                                                                                                                                                                                                                                                                                                            =          ?                 ^k�     �   =   @   ^      )            x_signed  := (others => '0');   )            z_signed  := (others => '0');�   <   >   ^      )            y_signed  := (others => '0');5�_�  |  ~          }   @       ����                                                                                                                                                                                                                                                                                                                            =          ?                 ^k�     �   ?   A   ^      ,            atan_signed  := (others => '0');5�_�  }            ~   7        ����                                                                                                                                                                                                                                                                                                                            @          7          V       ^k�     �   [   ]   ^          end process cordic_iter_proc;�   Z   \   ^            end if;�   Y   [   ^               end if;�   X   Z   ^                  end case;�   W   Y   ^      )                  state <= waitingEnable;�   V   X   ^                        dv_o  <= '0';�   U   W   ^      #               when waitingValid =>�   T   V   ^                        end if;�   S   U   ^      +                     state <= waitingValid;�   R   T   ^      $                     inv_o <= inv_i;�   Q   S   ^      "                     dv_o  <= '1';�   P   R   ^                              end if;�   O   Q   ^      =                           zip1 <= std_logic_vector(zis+cis);�   N   P   ^      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   M   O   ^      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   L   N   ^                              else�   K   M   ^      :                        zip1 <= std_logic_vector(zis-cis);�   J   L   ^      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   I   K   ^      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   H   J   ^      $                     if yis < 0 then�   G   I   ^      '                     cis := signed(ci);�   F   H   ^      '                     zis := signed(zi);�   E   G   ^      '                     xis := signed(xi);�   D   F   ^      '                     yis := signed(yi);�   C   E   ^      $                  if en_i = '1' then�   B   D   ^      $               when waitingEnable =>�   A   C   ^                  case state is�   @   B   ^               else�   ?   A   ^      +            atan_signed := (others => '0');�   >   @   ^      +            z_signed    := (others => '0');�   =   ?   ^      +            x_signed    := (others => '0');�   <   >   ^      +            y_signed    := (others => '0');�   ;   =   ^      +            m_dataZ     <= (others => '0');�   :   <   ^      +            m_dataY     <= (others => '0');�   9   ;   ^      +            m_dataX     <= (others => '0');�   8   :   ^      )            state       <= waitingEnable;�   7   9   ^                  s_inv       <= '0';�   6   8   ^                  s_ready     <= '0';�   5   7   ^               if rst = '0' then�   4   6   ^            if rising_edge(clk) then�   3   5   ^         begin�   2   4   ^      3      variable atan_signed : signed (N-1 downto 0);�   1   3   ^      3      variable z_signed    : signed (N-1 downto 0);�   0   2   ^      3      variable x_signed    : signed (N-1 downto 0);�   /   1   ^      3      variable y_signed    : signed (N-1 downto 0);�   .   0   ^      $   cordic_iter_proc:process (clk) is�   ,   .   ^      2   signal state:       stateType := waitingEnable;�   +   -   ^      4   type   stateType is (waitingValid,waitingEnable);�   '   )   ^                );�   &   (   ^      :--             zip1  : out std_logic_vector (N-1 downto 0)�   %   '   ^      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   $   &   ^      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   #   %   ^      %--             inv_o : out std_logic;�   "   $   ^      %--             dv_o  : out std_logic;�   !   #   ^      ;--             ci    : in  std_logic_vector (N-1 downto 0);�       "   ^      ;--             zi    : in  std_logic_vector (N-1 downto 0);�      !   ^      ;--             yi    : in  std_logic_vector (N-1 downto 0);�          ^      ;--             xi    : in  std_logic_vector (N-1 downto 0);�         ^      %--             inv_i : in  std_logic;�         ^      %--             en_i  : in  std_logic;�         ^      %--             rst   : in  std_logic;�         ^      %--             clk   : in  std_logic;�         ^      )          rst           : in  STD_LOGIC);�         ^      (          clk           : in  STD_LOGIC;�         ^      "          s_atan  : in  STD_LOGIC;�         ^      "          s_inv   : in  STD_LOGIC;�         ^      "          s_ready : out STD_LOGIC;�         ^      "          s_valid : in  STD_LOGIC;�         ^      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      "          m_ready : in  STD_LOGIC;�         ^      "          m_inv   : out STD_LOGIC;�         ^      "          m_valid : out STD_LOGIC;�         ^      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      ^      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      ^      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   ^            port(�      	   ^      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         ^      9             N     : natural := 16; --Ancho de la palabra�         ^            generic(�   6   8                      s_ready  <= '0';�   <   >          +            y_signed    := (others => '0');�   ;   =          '            m_dataZ <= (others => '0');�   ?   A          +            atan_signed := (others => '0');�   7   9                      s_inv <= '0';�   >   @          +            z_signed    := (others => '0');�   =   ?          +            x_signed    := (others => '0');�   :   <          '            m_dataY <= (others => '0');�   9   ;          '            m_dataX <= (others => '0');�   8   :          #            state <= waitingEnable;5�_�  ~  �             D       ����                                                                                                                                                                                                                                                                                                                            @          7          V       ^k�     �   C   E   ^      $                  if en_i = '1' then5�_�    �          �   D       ����                                                                                                                                                                                                                                                                                                                            @          7          V       ^k�     �   C   E   ^      +                  if s_validen_i = '1' then5�_�  �  �          �   D       ����                                                                                                                                                                                                                                                                                                                            @          7          V       ^l     �   C   E   ^      &                  if s_valid= '1' then5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l-     �   E   H   ^      '                     xis := signed(xi);   '                     zis := signed(zi);�   D   F   ^      '                     yis := signed(yi);5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l2     �   G   I   ^      '                     cis := signed(ci);5�_�  �  �          �   H        ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l5     �   G   I   ^      2                     atan_signedcis := signed(ci);5�_�  �  �          �   H        ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l5     �   G   I   ^      1                     atan_signedis := signed(ci);5�_�  �  �          �   H        ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l6     �   G   I   ^      0                     atan_signeds := signed(ci);5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            G          E                 ^l8     �   D   H   ^      .                     y_signedis := signed(yi);   .                     x_signedis := signed(xi);   .                     z_signedis := signed(zi);5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            E          G                 ^l:     �   E   H   ^      ,                     x_signed := signed(xi);   ,                     z_signed := signed(zi);�   D   F   ^      ,                     y_signed := signed(yi);5�_�  �  �          �   E        ����                                                                                                                                                                                                                                                                                                                            E          H          V       ^l=     �   [   ]   ^          end process cordic_iter_proc;�   Z   \   ^            end if;�   Y   [   ^               end if;�   X   Z   ^                  end case;�   W   Y   ^      )                  state <= waitingEnable;�   V   X   ^                        dv_o  <= '0';�   U   W   ^      #               when waitingValid =>�   T   V   ^                        end if;�   S   U   ^      +                     state <= waitingValid;�   R   T   ^      $                     inv_o <= inv_i;�   Q   S   ^      "                     dv_o  <= '1';�   P   R   ^                              end if;�   O   Q   ^      =                           zip1 <= std_logic_vector(zis+cis);�   N   P   ^      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   M   O   ^      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   L   N   ^                              else�   K   M   ^      :                        zip1 <= std_logic_vector(zis-cis);�   J   L   ^      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   I   K   ^      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   H   J   ^      $                     if yis < 0 then�   G   I   ^      /                     atan_signed := signed(ci);�   F   H   ^      /                     z_signed    := signed(zi);�   E   G   ^      /                     x_signed    := signed(xi);�   D   F   ^      /                     y_signed    := signed(yi);�   C   E   ^      '                  if s_valid = '1' then�   B   D   ^      $               when waitingEnable =>�   A   C   ^                  case state is�   @   B   ^               else�   ?   A   ^      +            atan_signed := (others => '0');�   >   @   ^      +            z_signed    := (others => '0');�   =   ?   ^      +            x_signed    := (others => '0');�   <   >   ^      +            y_signed    := (others => '0');�   ;   =   ^      +            m_dataZ     <= (others => '0');�   :   <   ^      +            m_dataY     <= (others => '0');�   9   ;   ^      +            m_dataX     <= (others => '0');�   8   :   ^      )            state       <= waitingEnable;�   7   9   ^                  s_inv       <= '0';�   6   8   ^                  s_ready     <= '0';�   5   7   ^               if rst = '0' then�   4   6   ^            if rising_edge(clk) then�   3   5   ^         begin�   2   4   ^      3      variable atan_signed : signed (N-1 downto 0);�   1   3   ^      3      variable z_signed    : signed (N-1 downto 0);�   0   2   ^      3      variable x_signed    : signed (N-1 downto 0);�   /   1   ^      3      variable y_signed    : signed (N-1 downto 0);�   .   0   ^      $   cordic_iter_proc:process (clk) is�   ,   .   ^      2   signal state:       stateType := waitingEnable;�   +   -   ^      4   type   stateType is (waitingValid,waitingEnable);�   '   )   ^                );�   &   (   ^      :--             zip1  : out std_logic_vector (N-1 downto 0)�   %   '   ^      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   $   &   ^      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   #   %   ^      %--             inv_o : out std_logic;�   "   $   ^      %--             dv_o  : out std_logic;�   !   #   ^      ;--             ci    : in  std_logic_vector (N-1 downto 0);�       "   ^      ;--             zi    : in  std_logic_vector (N-1 downto 0);�      !   ^      ;--             yi    : in  std_logic_vector (N-1 downto 0);�          ^      ;--             xi    : in  std_logic_vector (N-1 downto 0);�         ^      %--             inv_i : in  std_logic;�         ^      %--             en_i  : in  std_logic;�         ^      %--             rst   : in  std_logic;�         ^      %--             clk   : in  std_logic;�         ^      )          rst           : in  STD_LOGIC);�         ^      (          clk           : in  STD_LOGIC;�         ^      "          s_atan  : in  STD_LOGIC;�         ^      "          s_inv   : in  STD_LOGIC;�         ^      "          s_ready : out STD_LOGIC;�         ^      "          s_valid : in  STD_LOGIC;�         ^      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      "          m_ready : in  STD_LOGIC;�         ^      "          m_inv   : out STD_LOGIC;�         ^      "          m_valid : out STD_LOGIC;�         ^      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      ^      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      ^      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   ^            port(�      	   ^      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         ^      9             N     : natural := 16; --Ancho de la palabra�         ^            generic(�   D   F          /                     y_signed    := signed(yi);�   G   I          /                     atan_signed := signed(ci);�   F   H          /                     z_signed    := signed(zi);�   E   G          /                     x_signed    := signed(xi);5�_�  �  �          �   E   +    ����                                                                                                                                                                                                                                                                                                                            E   +       H   +          +    ^lX     �   E   I   ^      /                     x_signed    := signed(xi);   /                     z_signed    := signed(zi);   /                     atan_signed := signed(ci);�   D   F   ^      /                     y_signed    := signed(yi);5�_�  �  �          �   F   1    ����                                                                                                                                                                                                                                                                                                                            E   +       H   +          +    ^l^     �   E   G   ^      6                     x_signed    := signed(s_dataXxi);5�_�  �  �          �   G   1    ����                                                                                                                                                                                                                                                                                                                            E   +       H   +          +    ^l`     �   F   H   ^      6                     z_signed    := signed(s_dataXzi);5�_�  �  �          �   H   1    ����                                                                                                                                                                                                                                                                                                                            E   +       H   +          +    ^lg     �   G   I   ^      6                     atan_signed := signed(s_dataXci);5�_�  �  �          �   E   2    ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^lj     �   D   I   ^      6                     y_signed    := signed(s_dataXyi);   6                     x_signed    := signed(s_dataYxi);   6                     z_signed    := signed(s_dataZzi);   6                     atan_signed := signed(s_dataTci);5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^ll     �   G   I   ^      4                     atan_signed := signed(s_dataT);5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^lm     �   G   I   ^      3                     tan_signed := signed(s_dataT);5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^lm     �   G   I   ^      2                     tn_signed := signed(s_dataT);5�_�  �  �          �   @       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^lr     �   ?   A   ^      +            atan_signed := (others => '0');5�_�  �  �          �   @       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^lr     �   ?   A   ^      *            tan_signed := (others => '0');5�_�  �  �          �   @       ����                                                                                                                                                                                                                                                                                                                            H   2       E   3          3    ^ls     �   ?   A   ^      )            tn_signed := (others => '0');5�_�  �  �          �   7        ����                                                                                                                                                                                                                                                                                                                            7          @          V       ^lw     �   [   ]   ^          end process cordic_iter_proc;�   Z   \   ^            end if;�   Y   [   ^               end if;�   X   Z   ^                  end case;�   W   Y   ^      )                  state <= waitingEnable;�   V   X   ^                        dv_o  <= '0';�   U   W   ^      #               when waitingValid =>�   T   V   ^                        end if;�   S   U   ^      +                     state <= waitingValid;�   R   T   ^      $                     inv_o <= inv_i;�   Q   S   ^      "                     dv_o  <= '1';�   P   R   ^                              end if;�   O   Q   ^      =                           zip1 <= std_logic_vector(zis+cis);�   N   P   ^      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   M   O   ^      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   L   N   ^                              else�   K   M   ^      :                        zip1 <= std_logic_vector(zis-cis);�   J   L   ^      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   I   K   ^      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   H   J   ^      $                     if yis < 0 then�   G   I   ^      1                     t_signed := signed(s_dataT);�   F   H   ^      4                     z_signed    := signed(s_dataZ);�   E   G   ^      4                     x_signed    := signed(s_dataY);�   D   F   ^      4                     y_signed    := signed(s_dataX);�   C   E   ^      '                  if s_valid = '1' then�   B   D   ^      $               when waitingEnable =>�   A   C   ^                  case state is�   @   B   ^               else�   ?   A   ^      (            t_signed := (others => '0');�   >   @   ^      (            z_signed := (others => '0');�   =   ?   ^      (            x_signed := (others => '0');�   <   >   ^      (            y_signed := (others => '0');�   ;   =   ^      (            m_dataZ  <= (others => '0');�   :   <   ^      (            m_dataY  <= (others => '0');�   9   ;   ^      (            m_dataX  <= (others => '0');�   8   :   ^      &            state    <= waitingEnable;�   7   9   ^                  s_inv    <= '0';�   6   8   ^                  s_ready  <= '0';�   5   7   ^               if rst = '0' then�   4   6   ^            if rising_edge(clk) then�   3   5   ^         begin�   2   4   ^      3      variable atan_signed : signed (N-1 downto 0);�   1   3   ^      3      variable z_signed    : signed (N-1 downto 0);�   0   2   ^      3      variable x_signed    : signed (N-1 downto 0);�   /   1   ^      3      variable y_signed    : signed (N-1 downto 0);�   .   0   ^      $   cordic_iter_proc:process (clk) is�   ,   .   ^      2   signal state:       stateType := waitingEnable;�   +   -   ^      4   type   stateType is (waitingValid,waitingEnable);�   '   )   ^                );�   &   (   ^      :--             zip1  : out std_logic_vector (N-1 downto 0)�   %   '   ^      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   $   &   ^      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   #   %   ^      %--             inv_o : out std_logic;�   "   $   ^      %--             dv_o  : out std_logic;�   !   #   ^      ;--             ci    : in  std_logic_vector (N-1 downto 0);�       "   ^      ;--             zi    : in  std_logic_vector (N-1 downto 0);�      !   ^      ;--             yi    : in  std_logic_vector (N-1 downto 0);�          ^      ;--             xi    : in  std_logic_vector (N-1 downto 0);�         ^      %--             inv_i : in  std_logic;�         ^      %--             en_i  : in  std_logic;�         ^      %--             rst   : in  std_logic;�         ^      %--             clk   : in  std_logic;�         ^      )          rst           : in  STD_LOGIC);�         ^      (          clk           : in  STD_LOGIC;�         ^      "          s_atan  : in  STD_LOGIC;�         ^      "          s_inv   : in  STD_LOGIC;�         ^      "          s_ready : out STD_LOGIC;�         ^      "          s_valid : in  STD_LOGIC;�         ^      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      "          m_ready : in  STD_LOGIC;�         ^      "          m_inv   : out STD_LOGIC;�         ^      "          m_valid : out STD_LOGIC;�         ^      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      ^      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      ^      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   ^            port(�      	   ^      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         ^      9             N     : natural := 16; --Ancho de la palabra�         ^            generic(�   6   8                      s_ready     <= '0';�   <   >          +            y_signed    := (others => '0');�   ;   =          +            m_dataZ     <= (others => '0');�   ?   A          (            t_signed := (others => '0');�   7   9                      s_inv       <= '0';�   >   @          +            z_signed    := (others => '0');�   =   ?          +            x_signed    := (others => '0');�   :   <          +            m_dataY     <= (others => '0');�   9   ;          +            m_dataX     <= (others => '0');�   8   :          )            state       <= waitingEnable;5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            7          @          V       ^l|     �   2   4   ^      3      variable atan_signed : signed (N-1 downto 0);5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            7          @          V       ^l|     �   2   4   ^      2      variable tan_signed : signed (N-1 downto 0);5�_�  �  �          �   3       ����                                                                                                                                                                                                                                                                                                                            7          @          V       ^l}     �   2   4   ^      1      variable tn_signed : signed (N-1 downto 0);5�_�  �  �          �   0        ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^l~     �   [   ]   ^          end process cordic_iter_proc;�   Z   \   ^            end if;�   Y   [   ^               end if;�   X   Z   ^                  end case;�   W   Y   ^      )                  state <= waitingEnable;�   V   X   ^                        dv_o  <= '0';�   U   W   ^      #               when waitingValid =>�   T   V   ^                        end if;�   S   U   ^      +                     state <= waitingValid;�   R   T   ^      $                     inv_o <= inv_i;�   Q   S   ^      "                     dv_o  <= '1';�   P   R   ^                              end if;�   O   Q   ^      =                           zip1 <= std_logic_vector(zis+cis);�   N   P   ^      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   M   O   ^      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   L   N   ^                              else�   K   M   ^      :                        zip1 <= std_logic_vector(zis-cis);�   J   L   ^      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   I   K   ^      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   H   J   ^      $                     if yis < 0 then�   G   I   ^      1                     t_signed := signed(s_dataT);�   F   H   ^      4                     z_signed    := signed(s_dataZ);�   E   G   ^      4                     x_signed    := signed(s_dataY);�   D   F   ^      4                     y_signed    := signed(s_dataX);�   C   E   ^      '                  if s_valid = '1' then�   B   D   ^      $               when waitingEnable =>�   A   C   ^                  case state is�   @   B   ^               else�   ?   A   ^      (            t_signed := (others => '0');�   >   @   ^      (            z_signed := (others => '0');�   =   ?   ^      (            x_signed := (others => '0');�   <   >   ^      (            y_signed := (others => '0');�   ;   =   ^      (            m_dataZ  <= (others => '0');�   :   <   ^      (            m_dataY  <= (others => '0');�   9   ;   ^      (            m_dataX  <= (others => '0');�   8   :   ^      &            state    <= waitingEnable;�   7   9   ^                  s_inv    <= '0';�   6   8   ^                  s_ready  <= '0';�   5   7   ^               if rst = '0' then�   4   6   ^            if rising_edge(clk) then�   3   5   ^         begin�   2   4   ^      0      variable t_signed : signed (N-1 downto 0);�   1   3   ^      3      variable z_signed    : signed (N-1 downto 0);�   0   2   ^      3      variable x_signed    : signed (N-1 downto 0);�   /   1   ^      3      variable y_signed    : signed (N-1 downto 0);�   .   0   ^      $   cordic_iter_proc:process (clk) is�   ,   .   ^      2   signal state:       stateType := waitingEnable;�   +   -   ^      4   type   stateType is (waitingValid,waitingEnable);�   '   )   ^                );�   &   (   ^      :--             zip1  : out std_logic_vector (N-1 downto 0)�   %   '   ^      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   $   &   ^      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   #   %   ^      %--             inv_o : out std_logic;�   "   $   ^      %--             dv_o  : out std_logic;�   !   #   ^      ;--             ci    : in  std_logic_vector (N-1 downto 0);�       "   ^      ;--             zi    : in  std_logic_vector (N-1 downto 0);�      !   ^      ;--             yi    : in  std_logic_vector (N-1 downto 0);�          ^      ;--             xi    : in  std_logic_vector (N-1 downto 0);�         ^      %--             inv_i : in  std_logic;�         ^      %--             en_i  : in  std_logic;�         ^      %--             rst   : in  std_logic;�         ^      %--             clk   : in  std_logic;�         ^      )          rst           : in  STD_LOGIC);�         ^      (          clk           : in  STD_LOGIC;�         ^      "          s_atan  : in  STD_LOGIC;�         ^      "          s_inv   : in  STD_LOGIC;�         ^      "          s_ready : out STD_LOGIC;�         ^      "          s_valid : in  STD_LOGIC;�         ^      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      "          m_ready : in  STD_LOGIC;�         ^      "          m_inv   : out STD_LOGIC;�         ^      "          m_valid : out STD_LOGIC;�         ^      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      ^      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      ^      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   ^            port(�      	   ^      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         ^      9             N     : natural := 16; --Ancho de la palabra�         ^            generic(�   /   1          3      variable y_signed    : signed (N-1 downto 0);5�_�  �  �          �   0        ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^l�     �   [   ]   ^          end process cordic_iter_proc;�   Z   \   ^            end if;�   Y   [   ^               end if;�   X   Z   ^                  end case;�   W   Y   ^      )                  state <= waitingEnable;�   V   X   ^                        dv_o  <= '0';�   U   W   ^      #               when waitingValid =>�   T   V   ^                        end if;�   S   U   ^      +                     state <= waitingValid;�   R   T   ^      $                     inv_o <= inv_i;�   Q   S   ^      "                     dv_o  <= '1';�   P   R   ^                              end if;�   O   Q   ^      =                           zip1 <= std_logic_vector(zis+cis);�   N   P   ^      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   M   O   ^      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   L   N   ^                              else�   K   M   ^      :                        zip1 <= std_logic_vector(zis-cis);�   J   L   ^      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   I   K   ^      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   H   J   ^      $                     if yis < 0 then�   G   I   ^      1                     t_signed := signed(s_dataT);�   F   H   ^      4                     z_signed    := signed(s_dataZ);�   E   G   ^      4                     x_signed    := signed(s_dataY);�   D   F   ^      4                     y_signed    := signed(s_dataX);�   C   E   ^      '                  if s_valid = '1' then�   B   D   ^      $               when waitingEnable =>�   A   C   ^                  case state is�   @   B   ^               else�   ?   A   ^      (            t_signed := (others => '0');�   >   @   ^      (            z_signed := (others => '0');�   =   ?   ^      (            x_signed := (others => '0');�   <   >   ^      (            y_signed := (others => '0');�   ;   =   ^      (            m_dataZ  <= (others => '0');�   :   <   ^      (            m_dataY  <= (others => '0');�   9   ;   ^      (            m_dataX  <= (others => '0');�   8   :   ^      &            state    <= waitingEnable;�   7   9   ^                  s_inv    <= '0';�   6   8   ^                  s_ready  <= '0';�   5   7   ^               if rst = '0' then�   4   6   ^            if rising_edge(clk) then�   3   5   ^         begin�   2   4   ^      0      variable t_signed : signed (N-1 downto 0);�   1   3   ^      0      variable z_signed : signed (N-1 downto 0);�   0   2   ^      0      variable x_signed : signed (N-1 downto 0);�   /   1   ^      0      variable y_signed : signed (N-1 downto 0);�   .   0   ^      $   cordic_iter_proc:process (clk) is�   ,   .   ^      2   signal state:       stateType := waitingEnable;�   +   -   ^      4   type   stateType is (waitingValid,waitingEnable);�   '   )   ^                );�   &   (   ^      :--             zip1  : out std_logic_vector (N-1 downto 0)�   %   '   ^      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   $   &   ^      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   #   %   ^      %--             inv_o : out std_logic;�   "   $   ^      %--             dv_o  : out std_logic;�   !   #   ^      ;--             ci    : in  std_logic_vector (N-1 downto 0);�       "   ^      ;--             zi    : in  std_logic_vector (N-1 downto 0);�      !   ^      ;--             yi    : in  std_logic_vector (N-1 downto 0);�          ^      ;--             xi    : in  std_logic_vector (N-1 downto 0);�         ^      %--             inv_i : in  std_logic;�         ^      %--             en_i  : in  std_logic;�         ^      %--             rst   : in  std_logic;�         ^      %--             clk   : in  std_logic;�         ^      )          rst           : in  STD_LOGIC);�         ^      (          clk           : in  STD_LOGIC;�         ^      "          s_atan  : in  STD_LOGIC;�         ^      "          s_inv   : in  STD_LOGIC;�         ^      "          s_ready : out STD_LOGIC;�         ^      "          s_valid : in  STD_LOGIC;�         ^      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         ^      "          m_ready : in  STD_LOGIC;�         ^      "          m_inv   : out STD_LOGIC;�         ^      "          m_valid : out STD_LOGIC;�         ^      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      ^      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      ^      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   ^            port(�      	   ^      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         ^      9             N     : natural := 16; --Ancho de la palabra�         ^            generic(�   0   2          3      variable x_signed    : signed (N-1 downto 0);�   /   1          3      variable y_signed    : signed (N-1 downto 0);�   2   4          0      variable t_signed : signed (N-1 downto 0);�   1   3          3      variable z_signed    : signed (N-1 downto 0);5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^l�     �         ^    �         ^    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �         _      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �                8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            3          0          V       ^l�     �         ^    �         ^    5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �         _      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �         _      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �         _      8          s_dataU : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                            4          1          V       ^l�     �         _      8          s_dataE : in  STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �  �          �   F        ����                                                                                                                                                                                                                                                                                                                            I          F          V       ^l�     �   \   ^   _          end process cordic_iter_proc;�   [   ]   _            end if;�   Z   \   _               end if;�   Y   [   _                  end case;�   X   Z   _      )                  state <= waitingEnable;�   W   Y   _                        dv_o  <= '0';�   V   X   _      #               when waitingValid =>�   U   W   _                        end if;�   T   V   _      +                     state <= waitingValid;�   S   U   _      $                     inv_o <= inv_i;�   R   T   _      "                     dv_o  <= '1';�   Q   S   _                              end if;�   P   R   _      =                           zip1 <= std_logic_vector(zis+cis);�   O   Q   _      P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));�   N   P   _      P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));�   M   O   _                              else�   L   N   _      :                        zip1 <= std_logic_vector(zis-cis);�   K   M   _      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));�   J   L   _      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));�   I   K   _      $                     if yis < 0 then�   H   J   _      1                     t_signed := signed(s_dataT);�   G   I   _      1                     z_signed := signed(s_dataZ);�   F   H   _      1                     x_signed := signed(s_dataY);�   E   G   _      1                     y_signed := signed(s_dataX);�   D   F   _      '                  if s_valid = '1' then�   C   E   _      $               when waitingEnable =>�   B   D   _                  case state is�   A   C   _               else�   @   B   _      (            t_signed := (others => '0');�   ?   A   _      (            z_signed := (others => '0');�   >   @   _      (            x_signed := (others => '0');�   =   ?   _      (            y_signed := (others => '0');�   <   >   _      (            m_dataZ  <= (others => '0');�   ;   =   _      (            m_dataY  <= (others => '0');�   :   <   _      (            m_dataX  <= (others => '0');�   9   ;   _      &            state    <= waitingEnable;�   8   :   _                  s_inv    <= '0';�   7   9   _                  s_ready  <= '0';�   6   8   _               if rst = '0' then�   5   7   _            if rising_edge(clk) then�   4   6   _         begin�   3   5   _      0      variable t_signed : signed (N-1 downto 0);�   2   4   _      0      variable z_signed : signed (N-1 downto 0);�   1   3   _      0      variable x_signed : signed (N-1 downto 0);�   0   2   _      0      variable y_signed : signed (N-1 downto 0);�   /   1   _      $   cordic_iter_proc:process (clk) is�   -   /   _      2   signal state:       stateType := waitingEnable;�   ,   .   _      4   type   stateType is (waitingValid,waitingEnable);�   (   *   _                );�   '   )   _      :--             zip1  : out std_logic_vector (N-1 downto 0)�   &   (   _      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   %   '   _      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   $   &   _      %--             inv_o : out std_logic;�   #   %   _      %--             dv_o  : out std_logic;�   "   $   _      ;--             ci    : in  std_logic_vector (N-1 downto 0);�   !   #   _      ;--             zi    : in  std_logic_vector (N-1 downto 0);�       "   _      ;--             yi    : in  std_logic_vector (N-1 downto 0);�      !   _      ;--             xi    : in  std_logic_vector (N-1 downto 0);�          _      %--             inv_i : in  std_logic;�         _      %--             en_i  : in  std_logic;�         _      %--             rst   : in  std_logic;�         _      %--             clk   : in  std_logic;�         _      )          rst           : in  STD_LOGIC);�         _      (          clk           : in  STD_LOGIC;�         _      "          s_atan  : in  STD_LOGIC;�         _      "          s_inv   : in  STD_LOGIC;�         _      "          s_ready : out STD_LOGIC;�         _      "          s_valid : in  STD_LOGIC;�         _      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      "          m_ready : in  STD_LOGIC;�         _      "          m_inv   : out STD_LOGIC;�         _      "          m_valid : out STD_LOGIC;�         _      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      _      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      _      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   _            port(�      	   _      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         _      9             N     : natural := 16; --Ancho de la palabra�         _            generic(�   E   G          4                     y_signed    := signed(s_dataX);�   H   J          1                     t_signed := signed(s_dataT);�   G   I          4                     z_signed    := signed(s_dataZ);�   F   H          4                     x_signed    := signed(s_dataY);5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                            I          F          V       ^l�     �   I   K   _      $                     if yis < 0 then5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                            K          M                 ^l�     �   K   N   _      M                        yip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));   :                        zip1 <= std_logic_vector(zis-cis);�   J   L   _      M                        xip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));5�_�  �  �          �   K       ����                                                                                                                                                                                                                                                                                                                            K          M   "          "    ^l�     �   J   N   _      T                        m_dataXxip1 <= std_logic_vector(xis-shift_right(yis,SHIFT));   T                        m_dataXyip1 <= std_logic_vector(yis+shift_right(xis,SHIFT));   A                        m_dataXzip1 <= std_logic_vector(zis-cis);5�_�  �  �          �   L       ����                                                                                                                                                                                                                                                                                                                            K          M   "          "    ^l�     �   K   M   _      P                        m_dataX <= std_logic_vector(yis+shift_right(xis,SHIFT));5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                            K          M   "          "    ^l�     �   L   N   _      =                        m_dataX <= std_logic_vector(zis-cis);5�_�  �  �          �   K   4    ����                                                                                                                                                                                                                                                                                                                            K   4       M   4          4    ^m     �   K   N   _      P                        m_dataY <= std_logic_vector(yis+shift_right(xis,SHIFT));   =                        m_dataZ <= std_logic_vector(zis-cis);�   J   L   _      P                        m_dataX <= std_logic_vector(xis-shift_right(yis,SHIFT));5�_�  �  �          �   K   <    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m     �   J   N   _      X                        m_dataX <= std_logic_vector(x_signedxis-shift_right(yis,SHIFT));   X                        m_dataY <= std_logic_vector(x_signedyis+shift_right(xis,SHIFT));   E                        m_dataZ <= std_logic_vector(x_signedzis-cis);5�_�  �  �          �   L   4    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m     �   K   M   _      U                        m_dataY <= std_logic_vector(x_signed+shift_right(xis,SHIFT));5�_�  �  �          �   M   4    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m     �   L   N   _      B                        m_dataZ <= std_logic_vector(x_signed-cis);5�_�  �  �          �   K   I    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m     �   J   L   _      U                        m_dataX <= std_logic_vector(x_signed-shift_right(yis,SHIFT));5�_�  �  �          �   L   J    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m      �   K   M   _      U                        m_dataY <= std_logic_vector(y_signed+shift_right(xis,SHIFT));5�_�  �  �          �   L   Q    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m"     �   K   M   _      \                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signedis,SHIFT));5�_�  �  �          �   L   Q    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m"     �   K   M   _      [                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signeds,SHIFT));5�_�  �  �          �   M   =    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m$     �   L   N   _      B                        m_dataZ <= std_logic_vector(z_signed-cis);5�_�  �  �          �   M   E    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m&     �   L   N   _      J                        m_dataZ <= std_logic_vector(z_signed-t_signedcis);5�_�  �  �          �   M   E    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m&     �   L   N   _      I                        m_dataZ <= std_logic_vector(z_signed-t_signedis);5�_�  �  �          �   M   E    ����                                                                                                                                                                                                                                                                                                                            K   <       M   >          >    ^m'     �   L   N   _      H                        m_dataZ <= std_logic_vector(z_signed-t_signeds);5�_�  �  �          �   O        ����                                                                                                                                                                                                                                                                                                                            K          M          V       ^mZ     �   N   R   _    �   O   P   _    5�_�  �  �          �   O        ����                                                                                                                                                                                                                                                                                                                            O   !       Q   !       V   !    ^m]     �   P   R          G                        m_dataZ <= std_logic_vector(z_signed-t_signed);�   O   Q          Z                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signed,SHIFT));�   N   P          Z                        m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));5�_�  �  �          �   Q   ?    ����                                                                                                                                                                                                                                                                                                                            O   !       Q   !       V   !    ^ma     �   P   R   b      J                           m_dataZ <= std_logic_vector(z_signed-t_signed);5�_�  �  �          �   O   ?    ����                                                                                                                                                                                                                                                                                                                            O   !       Q   !       V   !    ^mf     �   N   P   b      ]                           m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));5�_�  �  �          �   P   ?    ����                                                                                                                                                                                                                                                                                                                            O   !       Q   !       V   !    ^mj     �   O   Q   b      ]                           m_dataY <= std_logic_vector(y_signed+shift_right(x_signed,SHIFT));5�_�  �  �          �   R        ����                                                                                                                                                                                                                                                                                                                            R   ?       T   =       V   ?    ^mm     �   Q   R          P                           xip1 <= std_logic_vector(xis+shift_right(yis,SHIFT));   P                           yip1 <= std_logic_vector(yis-shift_right(xis,SHIFT));   =                           zip1 <= std_logic_vector(zis+cis);5�_�  �  �          �   N        ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^ms     �   Q   S                                  end if;�   P   R          J                           m_dataZ <= std_logic_vector(z_signed+t_signed);�   O   Q          ]                           m_dataY <= std_logic_vector(y_signed-shift_right(x_signed,SHIFT));�   N   P          ]                           m_dataX <= std_logic_vector(x_signed+shift_right(y_signed,SHIFT));�   M   O                                  else5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^mx     �   R   T   _      "                     dv_o  <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   R   T   _      )                     m_validdv_o  <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   R   T   _      (                     m_validv_o  <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   R   T   _      '                     m_valid_o  <= '1';5�_�  �  �          �   S       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   R   T   _      &                     m_valido  <= '1';5�_�  �  �          �   T       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   S   U   _      $                     inv_o <= inv_i;5�_�  �  �          �   T       ����                                                                                                                                                                                                                                                                                                                            R          J          V       ^m�     �   S   U   _      $                     m_inv <= inv_i;5�_�  �  �          �   S        ����                                                                                                                                                                                                                                                                                                                            U          S          V       ^m�     �   \   ^   _          end process cordic_iter_proc;�   [   ]   _            end if;�   Z   \   _               end if;�   Y   [   _                  end case;�   X   Z   _      )                  state <= waitingEnable;�   W   Y   _                        dv_o  <= '0';�   V   X   _      #               when waitingValid =>�   U   W   _                        end if;�   T   V   _      -                     state   <= waitingValid;�   S   U   _      &                     m_inv   <= s_inv;�   R   T   _      $                     m_valid <= '1';�   Q   S   _                           end if;�   P   R   _      G                        m_dataZ <= std_logic_vector(z_signed+t_signed);�   O   Q   _      Z                        m_dataY <= std_logic_vector(y_signed-shift_right(x_signed,SHIFT));�   N   P   _      Z                        m_dataX <= std_logic_vector(x_signed+shift_right(y_signed,SHIFT));�   M   O   _                           else�   L   N   _      G                        m_dataZ <= std_logic_vector(z_signed-t_signed);�   K   M   _      Z                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signed,SHIFT));�   J   L   _      Z                        m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));�   I   K   _      )                     if y_signed < 0 then�   H   J   _      1                     t_signed := signed(s_dataT);�   G   I   _      1                     z_signed := signed(s_dataZ);�   F   H   _      1                     x_signed := signed(s_dataY);�   E   G   _      1                     y_signed := signed(s_dataX);�   D   F   _      '                  if s_valid = '1' then�   C   E   _      $               when waitingEnable =>�   B   D   _                  case state is�   A   C   _               else�   @   B   _      (            t_signed := (others => '0');�   ?   A   _      (            z_signed := (others => '0');�   >   @   _      (            x_signed := (others => '0');�   =   ?   _      (            y_signed := (others => '0');�   <   >   _      (            m_dataZ  <= (others => '0');�   ;   =   _      (            m_dataY  <= (others => '0');�   :   <   _      (            m_dataX  <= (others => '0');�   9   ;   _      &            state    <= waitingEnable;�   8   :   _                  s_inv    <= '0';�   7   9   _                  s_ready  <= '0';�   6   8   _               if rst = '0' then�   5   7   _            if rising_edge(clk) then�   4   6   _         begin�   3   5   _      0      variable t_signed : signed (N-1 downto 0);�   2   4   _      0      variable z_signed : signed (N-1 downto 0);�   1   3   _      0      variable x_signed : signed (N-1 downto 0);�   0   2   _      0      variable y_signed : signed (N-1 downto 0);�   /   1   _      $   cordic_iter_proc:process (clk) is�   -   /   _      2   signal state:       stateType := waitingEnable;�   ,   .   _      4   type   stateType is (waitingValid,waitingEnable);�   (   *   _                );�   '   )   _      :--             zip1  : out std_logic_vector (N-1 downto 0)�   &   (   _      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   %   '   _      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   $   &   _      %--             inv_o : out std_logic;�   #   %   _      %--             dv_o  : out std_logic;�   "   $   _      ;--             ci    : in  std_logic_vector (N-1 downto 0);�   !   #   _      ;--             zi    : in  std_logic_vector (N-1 downto 0);�       "   _      ;--             yi    : in  std_logic_vector (N-1 downto 0);�      !   _      ;--             xi    : in  std_logic_vector (N-1 downto 0);�          _      %--             inv_i : in  std_logic;�         _      %--             en_i  : in  std_logic;�         _      %--             rst   : in  std_logic;�         _      %--             clk   : in  std_logic;�         _      )          rst           : in  STD_LOGIC);�         _      (          clk           : in  STD_LOGIC;�         _      "          s_atan  : in  STD_LOGIC;�         _      "          s_inv   : in  STD_LOGIC;�         _      "          s_ready : out STD_LOGIC;�         _      "          s_valid : in  STD_LOGIC;�         _      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      "          m_ready : in  STD_LOGIC;�         _      "          m_inv   : out STD_LOGIC;�         _      "          m_valid : out STD_LOGIC;�         _      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      _      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      _      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   _            port(�      	   _      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         _      9             N     : natural := 16; --Ancho de la palabra�         _            generic(�   R   T          %                     m_valid  <= '1';�   T   V          +                     state <= waitingValid;�   S   U          $                     m_inv <= s_inv;5�_�  �  �          �   X       ����                                                                                                                                                                                                                                                                                                                            U          S          V       ^m�     �   W   Y   _                        dv_o  <= '0';5�_�  �  �          �   X        ����                                                                                                                                                                                                                                                                                                                            Y          X          V       ^m�   0 �   \   ^   _          end process cordic_iter_proc;�   [   ]   _            end if;�   Z   \   _               end if;�   Y   [   _                  end case;�   X   Z   _      +                  state   <= waitingEnable;�   W   Y   _      !                  m_valid <= '0';�   V   X   _      #               when waitingValid =>�   U   W   _                        end if;�   T   V   _      -                     state   <= waitingValid;�   S   U   _      &                     m_inv   <= s_inv;�   R   T   _      $                     m_valid <= '1';�   Q   S   _                           end if;�   P   R   _      G                        m_dataZ <= std_logic_vector(z_signed+t_signed);�   O   Q   _      Z                        m_dataY <= std_logic_vector(y_signed-shift_right(x_signed,SHIFT));�   N   P   _      Z                        m_dataX <= std_logic_vector(x_signed+shift_right(y_signed,SHIFT));�   M   O   _                           else�   L   N   _      G                        m_dataZ <= std_logic_vector(z_signed-t_signed);�   K   M   _      Z                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signed,SHIFT));�   J   L   _      Z                        m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));�   I   K   _      )                     if y_signed < 0 then�   H   J   _      1                     t_signed := signed(s_dataT);�   G   I   _      1                     z_signed := signed(s_dataZ);�   F   H   _      1                     x_signed := signed(s_dataY);�   E   G   _      1                     y_signed := signed(s_dataX);�   D   F   _      '                  if s_valid = '1' then�   C   E   _      $               when waitingEnable =>�   B   D   _                  case state is�   A   C   _               else�   @   B   _      (            t_signed := (others => '0');�   ?   A   _      (            z_signed := (others => '0');�   >   @   _      (            x_signed := (others => '0');�   =   ?   _      (            y_signed := (others => '0');�   <   >   _      (            m_dataZ  <= (others => '0');�   ;   =   _      (            m_dataY  <= (others => '0');�   :   <   _      (            m_dataX  <= (others => '0');�   9   ;   _      &            state    <= waitingEnable;�   8   :   _                  s_inv    <= '0';�   7   9   _                  s_ready  <= '0';�   6   8   _               if rst = '0' then�   5   7   _            if rising_edge(clk) then�   4   6   _         begin�   3   5   _      0      variable t_signed : signed (N-1 downto 0);�   2   4   _      0      variable z_signed : signed (N-1 downto 0);�   1   3   _      0      variable x_signed : signed (N-1 downto 0);�   0   2   _      0      variable y_signed : signed (N-1 downto 0);�   /   1   _      $   cordic_iter_proc:process (clk) is�   -   /   _      2   signal state:       stateType := waitingEnable;�   ,   .   _      4   type   stateType is (waitingValid,waitingEnable);�   (   *   _                );�   '   )   _      :--             zip1  : out std_logic_vector (N-1 downto 0)�   &   (   _      ;--             yip1  : out std_logic_vector (N-1 downto 0);�   %   '   _      ;--             xip1  : out std_logic_vector (N-1 downto 0);�   $   &   _      %--             inv_o : out std_logic;�   #   %   _      %--             dv_o  : out std_logic;�   "   $   _      ;--             ci    : in  std_logic_vector (N-1 downto 0);�   !   #   _      ;--             zi    : in  std_logic_vector (N-1 downto 0);�       "   _      ;--             yi    : in  std_logic_vector (N-1 downto 0);�      !   _      ;--             xi    : in  std_logic_vector (N-1 downto 0);�          _      %--             inv_i : in  std_logic;�         _      %--             en_i  : in  std_logic;�         _      %--             rst   : in  std_logic;�         _      %--             clk   : in  std_logic;�         _      )          rst           : in  STD_LOGIC);�         _      (          clk           : in  STD_LOGIC;�         _      "          s_atan  : in  STD_LOGIC;�         _      "          s_inv   : in  STD_LOGIC;�         _      "          s_ready : out STD_LOGIC;�         _      "          s_valid : in  STD_LOGIC;�         _      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         _      "          m_ready : in  STD_LOGIC;�         _      "          m_inv   : out STD_LOGIC;�         _      "          m_valid : out STD_LOGIC;�         _      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      _      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�   	      _      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�      
   _            port(�      	   _      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �         _      9             N     : natural := 16; --Ancho de la palabra�         _            generic(�   W   Y          "                  m_valid  <= '0';�   X   Z          )                  state <= waitingEnable;5�_�  �  �          �      
    ����                                                                                                                                                                                                                                                                                                                            )   
          
       V   
    ^u!   1 �                %--             clk   : in  std_logic;   %--             rst   : in  std_logic;   %--             en_i  : in  std_logic;   %--             inv_i : in  std_logic;   ;--             xi    : in  std_logic_vector (N-1 downto 0);   ;--             yi    : in  std_logic_vector (N-1 downto 0);   ;--             zi    : in  std_logic_vector (N-1 downto 0);   ;--             ci    : in  std_logic_vector (N-1 downto 0);   %--             dv_o  : out std_logic;   %--             inv_o : out std_logic;   ;--             xip1  : out std_logic_vector (N-1 downto 0);   ;--             yip1  : out std_logic_vector (N-1 downto 0);   :--             zip1  : out std_logic_vector (N-1 downto 0)             );5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^un   2 �                "          s_atan  : in  STD_LOGIC;5�_�  �  �  �      �   *       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^u�     �   )   +   P                  s_inv    <= '0';5�_�  �  �          �   *       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^u�   3 �   )   +   P                  m_inv    <= '0';5�_�  �  �          �   7       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^�@     �   6   8   P      1                     y_signed := signed(s_dataX);5�_�  �  �          �   8       ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^�A   4 �   7   9   P      1                     x_signed := signed(s_dataY);5�_�  �  �          �   E        ����                                                                                                                                                                                                                                                                                                                            E          E          V       ^��     �   D   E          &                     m_inv   <= s_inv;5�_�  �  �          �   D       ����                                                                                                                                                                                                                                                                                                                            E          E          V       ^��     �   C   E   O    �   D   E   O    5�_�  �  �          �   E       ����                                                                                                                                                                                                                                                                                                                            F          F          V       ^��     �   E   G   Q                           �   E   G   P    5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            G          G          V       ^��     �   E   G   Q                           if(m_ready5�_�  �  �          �   F       ����                                                                                                                                                                                                                                                                                                                            G          G          V       ^��     �   E   G   Q      %                     if(m_ready = '1'5�_�  �  �          �   F   %    ����                                                                                                                                                                                                                                                                                                                            G          G          V       ^��     �   E   G   Q      %                     if m_ready = '1'5�_�  �  �          �   G   )    ����                                                                                                                                                                                                                                                                                                                            G          G          V       ^��     �   F   H   Q    �   G   H   Q    5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            H          H          V       ^��     �   F   H          -                     state   <= waitingValid;5�_�  �  �          �   G   *    ����                                                                                                                                                                                                                                                                                                                            H          H          V       ^��     �   F   H   R      0                        state   <= waitingValid;5�_�  �  �          �   G   /    ����                                                                                                                                                                                                                                                                                                                            H          H          V       ^��     �   G   I   S                              �   G   I   R    5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            I          I          V       ^��     �   H   J          -                     state   <= waitingValid;5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                            I          I          V       ^��     �   I   K   S    �   J   K   S    5�_�  �  �          �   J       ����                                                                                                                                                                                                                                                                                                                            I          I          V       ^��     �   I   K                            end if;5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            I          I          V       ^��     �   H   J   T    �   I   J   T    5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^��     �   H   J          !                  m_valid <= '0';5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�l     �   H   J   U      '                        m_valid <= '0';5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�m     �   H   J   U      '                        s_valid <= '0';5�_�  �  �  �      �   )       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^��     �   (   *   U                  s_ready  <= '0';5�_�  �  �          �   G       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^��     �   F   H   U    �   G   H   U    5�_�  �  �          �   G   $    ����                                                                                                                                                                                                                                                                                                                            K          K          V       ^��     �   F   H   V      '                        s_ready <= '0';5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            K          K          V       ^��     �   G   H          1                        state   <= waitingEnable;5�_�  �  �  �      �   5       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�I     �   4   6   U      $               when waitingEnable =>5�_�  �  �          �   J   *    ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�R     �   I   K   U      0                        state   <= waitingValid;5�_�  �  �          �   M       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�U     �   L   N   U      #               when waitingValid =>5�_�  �  �          �   O   $    ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�W     �   N   P   U      +                  state   <= waitingEnable;5�_�  �  �          �      ,    ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�b     �         U      4   type   stateType is (waitingValid,waitingEnable);5�_�  �  �          �      +    ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�e     �          U      2   signal state:       stateType := waitingEnable;5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�k     �   *   ,   U      &            state    <= waitingEnable;5�_�  �  �          �   +        ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�l     �   *   ,   U      !            state    <= waitingV;5�_�  �  �          �   *       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^�z     �   )   +   U    �   *   +   U    5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            K          K          V       ^�{     �   *   ,   V                  m_inv    <= '0';5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            K          K          V       ^�~     �   *   ,   V                  m_valid    <= '0';5�_�  �  �          �   +       ����                                                                                                                                                                                                                                                                                                                            K          K          V       ^�~     �   *   ,   V                  m_valid   <= '0';5�_�  �  �          �   P        ����                                                                                                                                                                                                                                                                                                                            G          L          V       ^��     �   O   V   V    �   P   Q   V    5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            G          L          V       ^��     �   Q   S   \    �   R   S   \    5�_�  �  �          �   R   *    ����                                                                                                                                                                                                                                                                                                                            R   *       R   .       v   .    ^��     �   Q   S   ]      0                        state   <= waitingReady;5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            R   *       R   .       v   .    ^��     �   H   J   ]    �   I   J   ]    5�_�  �  �          �   I       ����                                                                                                                                                                                                                                                                                                                            S   *       S   .       v   .    ^��     �   H   I          0                        state   <= waitingValid;5�_�  �  �          �   G   #    ����                                                                                                                                                                                                                                                                                                                            R   *       R   .       v   .    ^��     �   F   H   ]      *                     if m_ready = '1' then5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            R   *       R   .       v   .    ^��     �   G   H          '                        s_ready <= '1';5�_�  �  �          �   H       ����                                                                                                                                                                                                                                                                                                                            Q   *       Q   .       v   .    ^��     �   G   H                               else5�_�  �  �          �   Q        ����                                                                                                                                                                                                                                                                                                                            Q          S          V       ^��     �   P   Q                               else   '                        s_ready <= '0';   0                        state   <= waitingReady;5�_�  �  �          �   R       ����                                                                                                                                                                                                                                                                                                                            Q          Q          V       ^��     �   Q   R          *                  state   <= waitingValid;5�_�  �             �   N       ����                                                                                                                                                                                                                                                                                                                            Q          N          V       ^��   7 �   P   R                               end if;�   O   Q          0                        state   <= waitingValid;�   N   P          '                        s_ready <= '1';�   M   O          *                     if m_ready = '1' then5�_�  �    �          K       ����                                                                                                                                                                                                                                                                                                                            Q          N          V       ^��     �   K   M   X                        �   K   M   W    5�_�                  K       ����                                                                                                                                                                                                                                                                                                                            R          O          V       ^��     �   J   M   Y                           �   J   L   X    5�_�                 L        ����                                                                                                                                                                                                                                                                                                                            L          L          V       ^��     �   K   M   Y    �   L   M   Y    �   K   L                               k5�_�                 L   !    ����                                                                                                                                                                                                                                                                                                                            L           L   #       V       ^��     �   K   M   Z      $                     m_valid <= '1';5�_�                 N       ����                                                                                                                                                                                                                                                                                                                            L           L   #       V       ^��   8 �   M   N                            kk5�_�                 O        ����                                                                                                                                                                                                                                                                                                                            O          O          V       ^��     �   N   O          !                  m_valid <= '0';5�_�                 P       ����                                                                                                                                                                                                                                                                                                                            O          O          V       ^��     �   O   Q   X    �   P   Q   X    5�_�                 P       ����                                                                                                                                                                                                                                                                                                                            O          O          V       ^��   < �   O   Q          !                  m_valid <= '0';5�_�    	             6        ����                                                                                                                                                                                                                                                                                                                            P          P          V       ^��     �   6   7   Y    �   5   6   Y      #               when waitingValid =>5�_�    
          	   6       ����                                                                                                                                                                                                                                                                                                                            P          P          V       ^��     �   5   7   Z      "               when waitingPipe =>5�_�  	            
   6       ����                                                                                                                                                                                                                                                                                                                            Q          Q          V       ^��     �   6   7   Z       5�_�  
               7        ����                                                                                                                                                                                                                                                                                                                            Q          Q          V       ^��     �   6   8   [      .                  bitCounter := bitCounter +1;5�_�                 7   -    ����                                                                                                                                                                                                                                                                                                                            S          S          V       ^��     �   7   8   [                        �   7   9   \      (                  if bitCounter = N then   +                     state := waitingValid;5�_�                 9   *    ����                                                                                                                                                                                                                                                                                                                            T          T          V       ^�#     �   9   :   ]                           �   9   ;   ^                        end if;5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            U          U          V       ^�-     �   4   5   ^    �   3   4   ^      .                  bitCounter := bitCounter +1;5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            U          U          V       ^�.     �   3   5          (            bitCounter := bitCounter +1;5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�0     �   3   5   _                  bitCounter := - +1;5�_�                 4       ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�3   : �   3   5   _                  bitCounter := 0;5�_�                 8   ,    ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�L   ; �   7   9   _      /                  bitCounter := bitCounter + 1;5�_�                 ,       ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�T     �   +   -   _      $            state    <= waitingPipe;5�_�                    1    ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�Y     �         _      @   type   stateType is (waitingValid,waitingReady, waitingPipe);5�_�                    +    ����                                                                                                                                                                                                                                                                                                                            4          4          v       ^�`     �          _      0   signal state:       stateType := waitingPipe;5�_�                 9   "    ����                                                                                                                                                                                                                                                                                                                            7   !       ;          V   "    ^��     �   8   :   _      ,                  if bitCounter = SHIFT then5�_�                   7        ����                                                                                                                                                                                                                                                                                                                            7   !       7          V   "    ^��     �   6   <        5�_�  �             �   K       ����                                                                                                                                                                                                                                                                                                                            R          O          V       ^��     �   K   L   W    �   K   L   W      T            s_validW(0)   <= '0';                           --y ya no tengo mas nada5�_�  �  �  �  �  �   J       ����                                                                                                                                                                                                                                                                                                                            D          E          V       ^��   5 �   I   K        5�_�  �      �      �   D        ����                                                                                                                                                                                                                                                                                                                            D          E          V       ^��   6 �   D   F          $                     m_valid <= '1';�   C   E          &                     m_inv   <= s_inv;�         T            generic(�         T      9             N     : natural := 16; --Ancho de la palabra�      	   T      v             SHIFT : natural := 1); -- en el for generate va tomando valores en funcion de la posicion en el pipeline �      
   T            port(�   	      T      8          m_dataX : out STD_LOGIC_VECTOR (N-1 downto 0);�   
      T      8          m_dataY : out STD_LOGIC_VECTOR (N-1 downto 0);�         T      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);�         T      "          m_valid : out STD_LOGIC;�         T      "          m_inv   : out STD_LOGIC;�         T      "          m_ready : in  STD_LOGIC;�         T      8          s_dataX : in  STD_LOGIC_VECTOR (N-1 downto 0);�         T      8          s_dataY : in  STD_LOGIC_VECTOR (N-1 downto 0);�         T      8          s_dataZ : in  STD_LOGIC_VECTOR (N-1 downto 0);�         T      8          s_dataT : in  STD_LOGIC_VECTOR (N-1 downto 0);�         T      "          s_valid : in  STD_LOGIC;�         T      "          s_ready : out STD_LOGIC;�         T      "          s_inv   : in  STD_LOGIC;�         T      (          clk           : in  STD_LOGIC;�         T      )          rst           : in  STD_LOGIC);�         T      4   type   stateType is (waitingValid,waitingEnable);�          T      2   signal state:       stateType := waitingEnable;�       "   T      $   cordic_iter_proc:process (clk) is�   !   #   T      0      variable y_signed : signed (N-1 downto 0);�   "   $   T      0      variable x_signed : signed (N-1 downto 0);�   #   %   T      0      variable z_signed : signed (N-1 downto 0);�   $   &   T      0      variable t_signed : signed (N-1 downto 0);�   %   '   T         begin�   &   (   T            if rising_edge(clk) then�   '   )   T               if rst = '0' then�   (   *   T                  s_ready  <= '1';�   )   +   T                  m_inv    <= '0';�   *   ,   T      &            state    <= waitingEnable;�   +   -   T      (            m_dataX  <= (others => '0');�   ,   .   T      (            m_dataY  <= (others => '0');�   -   /   T      (            m_dataZ  <= (others => '0');�   .   0   T      (            y_signed := (others => '0');�   /   1   T      (            x_signed := (others => '0');�   0   2   T      (            z_signed := (others => '0');�   1   3   T      (            t_signed := (others => '0');�   2   4   T               else�   3   5   T                  case state is�   4   6   T      $               when waitingEnable =>�   5   7   T      '                  if s_valid = '1' then�   6   8   T      1                     x_signed := signed(s_dataX);�   7   9   T      1                     y_signed := signed(s_dataY);�   8   :   T      1                     z_signed := signed(s_dataZ);�   9   ;   T      1                     t_signed := signed(s_dataT);�   :   <   T      )                     if y_signed < 0 then�   ;   =   T      Z                        m_dataX <= std_logic_vector(x_signed-shift_right(y_signed,SHIFT));�   <   >   T      Z                        m_dataY <= std_logic_vector(y_signed+shift_right(x_signed,SHIFT));�   =   ?   T      G                        m_dataZ <= std_logic_vector(z_signed-t_signed);�   >   @   T                           else�   ?   A   T      Z                        m_dataX <= std_logic_vector(x_signed+shift_right(y_signed,SHIFT));�   @   B   T      Z                        m_dataY <= std_logic_vector(y_signed-shift_right(x_signed,SHIFT));�   A   C   T      G                        m_dataZ <= std_logic_vector(z_signed+t_signed);�   B   D   T                           end if;�   C   E   T      &                     m_inv   <= s_inv;�   D   F   T      $                     m_valid <= '1';�   E   G   T      *                     if m_ready = '1' then�   F   H   T      '                        s_ready <= '1';�   G   I   T                           else�   H   J   T      '                        s_ready <= '0';�   I   K   T                           end if;�   J   L   T                        end if;�   K   M   T      #               when waitingValid =>�   L   N   T      !                  m_valid <= '0';�   M   O   T      +                  state   <= waitingEnable;�   N   P   T                  end case;�   O   Q   T               end if;�   P   R   T            end if;�   Q   S   T          end process cordic_iter_proc;5�_�  �          �  �   D       ����                                                                                                                                                                                                                                                                                                                            E          D          V       ^��     �   C   F   T      &eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   $eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee5�_�  �          �  �   H       ����                                                                                                                                                                                                                                                                                                                            H          H          V       ^��     �   G   J        5�_�  �          �  �   (       ����                                                                                                                                                                                                                                                                                                                            J          J          V       ^��     �   '   )   U               if rst = '0' the15�_�  �  �      �  �           ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^uq     �         P    �         P      8          m_dataZ : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                               
          
       V   
    ^ut     �         Q      8          m_dataT : out STD_LOGIC_VECTOR (N-1 downto 0);5�_�  d          f  e      
    ����                                                                                                                                                                                                                                                                                                                            0   (       3   )          )    ^k�     �         ^                 : out STD_LOGIC;5�_�               ,        ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�r     �   +   -        5�_�                   ,   	    ����                                                                                                                                                                                                                                                                                                                            )          )          V       ^�s     �   ,   -   H       5�_�   �           �   �   !       ����                                                                                                                                                                                                                                                                                                                            &          !          V       ^�#     �       '   <      eeeeeeeeeeeeeeeeeeeeeeeee   #eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   #eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   #eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   #eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee   eeeeeeeeeeeeeeeeeeeee5�_�   j           l   k   )        ����                                                                                                                                                                                                                                                                                                                            )           )           V        ^�Y     �   (   .        5�_�   <   >       @   =   (       ����                                                                                                                                                                                                                                                                                                                            -          -          v       ^�~     �   (   )   4    �   '   (   4      !                     dv_o <= '1';5�_�   =   ?           >   (       ����                                                                                                                                                                                                                                                                                                                            -          -          v       ^��     �   '   )   5      !                     dv_o <= '-';5�_�   >               ?   +       ����                                                                                                                                                                                                                                                                                                                            .          .          v       ^��     �   +   ,   5                           �   +   -   6                        else5�_�   2           4   3   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v       ^�&     �   +   -   3      #               when waitingVali =>5�_�   %           '   &   %       ����                                                                                                                                                                                                                                                                                                                            $          $          v       ^��     �   %   &   .    �   $   &   .               else: stateType5�_�                    &       ����                                                                                                                                                                                                                                                                                                                            #          #          v       ^�?     �   %   '   (      !   end process cordic_'iter_proc;5��