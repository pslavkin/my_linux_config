Vim�UnDo� �1"���V���e^��='M<I����:)h��   L   +architecture Behavioral of slice_8from47 is      '   b   t          t   t    ^2]�    _�       c           b      1    ����                                                                                                                                                                                                                                                                                                                                                             ^2SS     �         L      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (31 downto 0);5�_�   b   d           c      2    ����                                                                                                                                                                                                                                                                                                                                                             ^2SU     �         L      >           s_axis_tdata  : in  STD_LOGIC_VECTOR (48 downto 0);5�_�   c   e           d      &    ����                                                                                                                                                                                                                                                                                                                                                             ^2SY     �         L      +architecture Behavioral of slice_8from32 is5�_�   d   f           e   /   &    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2Sw     �   .   0   L      T                     m_axis_tdata  <= s_axis_tdata(30) & s_axis_tdata(30 downto 24);5�_�   e   g           f   /   3    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2Sz     �   .   0   L      A                     m_axis_tdata  <= s_axis_tdata(30 downto 24);5�_�   f   h           g   /   =    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   .   0   L      A                     m_axis_tdata  <= s_axis_tdata(45 downto 24);5�_�   g   i           h   8   6    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   7   9   L      D                        m_axis_tdata  <= s_axis_tdata(23 downto 16);5�_�   h   j           i   8   @    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   7   9   L      D                        m_axis_tdata  <= s_axis_tdata(37 downto 16);5�_�   i   k           j   :   6    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      V                        m_axis_tdata  <= s_axis_tdata(14) & s_axis_tdata(14 downto 8);5�_�   j   l           k   :   I    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      V                        m_axis_tdata  <= s_axis_tdata(21) & s_axis_tdata(14 downto 8);5�_�   k   m           l   :   S    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      V                        m_axis_tdata  <= s_axis_tdata(21) & s_axis_tdata(21 downto 8);5�_�   l   n           m   :   )    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      W                        m_axis_tdata  <= s_axis_tdata(21) & s_axis_tdata(21 downto 14);5�_�   m   o           n   :   )    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      F                        m_axis_tdata  <= & s_axis_tdata(21 downto 14);5�_�   n   p           o   :   )    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   9   ;   L      E                        m_axis_tdata  <=  s_axis_tdata(21 downto 14);5�_�   o   q           p   <   6    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�     �   ;   =   L      B                        m_axis_tdata  <= s_axis_tdata(7 downto 0);5�_�   p   r           q   <   @    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2S�    �   ;   =   L      C                        m_axis_tdata  <= s_axis_tdata(13 downto 0);5�_�   q   s           r          ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2T%     �         L      entity slice_8from32 is5�_�   r   t           s          ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2T+    �         L      end slice_8from32;5�_�   s               t      '    ����                                                                                                                                                                                                                                                                                                                            /   &       /   8       v   8    ^2]�    �         L      +architecture Behavioral of slice_8from47 is5��